magic
tech scmos
timestamp 1732045399
<< nwell >>
rect -336 -377 -304 -251
rect -284 -377 -252 -251
rect -232 -315 -200 -251
rect -180 -315 -148 -251
rect -132 -361 -68 -297
rect 1571 -391 1603 -265
rect 1623 -391 1655 -265
rect 1675 -329 1707 -265
rect 1727 -329 1759 -265
rect 1775 -375 1839 -311
rect 144 -475 168 -455
rect 174 -475 230 -455
rect -339 -604 -307 -478
rect -287 -604 -255 -478
rect -235 -542 -203 -478
rect -183 -542 -151 -478
rect -135 -588 -71 -524
rect 144 -525 168 -505
rect 957 -545 981 -525
rect 987 -545 1043 -525
rect 145 -596 169 -576
rect 175 -596 231 -576
rect 957 -595 981 -575
rect 145 -646 169 -626
rect 625 -654 667 -620
rect 709 -659 733 -635
rect 778 -659 812 -623
rect 1563 -633 1595 -507
rect 1615 -633 1647 -507
rect 1667 -571 1699 -507
rect 1719 -571 1751 -507
rect 1767 -617 1831 -553
rect 819 -660 843 -636
rect 967 -669 991 -649
rect 997 -669 1053 -649
rect -342 -833 -310 -707
rect -290 -833 -258 -707
rect -238 -771 -206 -707
rect -186 -771 -154 -707
rect 145 -717 169 -697
rect 175 -717 231 -697
rect 489 -745 541 -697
rect 547 -743 577 -703
rect 967 -719 991 -699
rect -138 -817 -74 -753
rect 145 -767 169 -747
rect 601 -779 635 -743
rect 642 -780 666 -756
rect 145 -837 169 -817
rect 175 -837 231 -817
rect 488 -845 528 -811
rect 871 -823 895 -803
rect 901 -823 957 -803
rect 565 -850 589 -826
rect 145 -887 169 -867
rect 640 -887 674 -851
rect 681 -888 705 -864
rect 871 -873 895 -853
rect 1564 -869 1596 -743
rect 1616 -869 1648 -743
rect 1668 -807 1700 -743
rect 1720 -807 1752 -743
rect 1768 -853 1832 -789
rect -342 -1049 -310 -923
rect -290 -1049 -258 -923
rect -238 -987 -206 -923
rect -186 -987 -154 -923
rect -138 -1033 -74 -969
rect 846 -1015 886 -981
rect 924 -1020 948 -996
rect 165 -1088 205 -1054
rect 243 -1093 267 -1069
rect 1000 -1082 1034 -1046
rect 1041 -1083 1065 -1059
rect 850 -1122 890 -1088
rect 928 -1127 952 -1103
rect 1315 -1109 1339 -1089
rect 1345 -1109 1401 -1089
rect 1564 -1102 1596 -976
rect 1616 -1102 1648 -976
rect 1668 -1040 1700 -976
rect 1720 -1040 1752 -976
rect 1768 -1086 1832 -1022
rect -343 -1264 -311 -1138
rect -291 -1264 -259 -1138
rect -239 -1202 -207 -1138
rect -187 -1202 -155 -1138
rect 166 -1175 206 -1141
rect 243 -1180 267 -1156
rect 1088 -1161 1122 -1125
rect 1129 -1162 1153 -1138
rect 1315 -1159 1339 -1139
rect -139 -1248 -75 -1184
rect 168 -1263 208 -1229
rect 850 -1231 890 -1197
rect 928 -1236 952 -1212
rect 246 -1268 270 -1244
rect 1000 -1251 1034 -1215
rect 1041 -1252 1065 -1228
rect 168 -1349 208 -1315
rect 1559 -1328 1591 -1202
rect 1611 -1328 1643 -1202
rect 1663 -1266 1695 -1202
rect 1715 -1266 1747 -1202
rect 1763 -1312 1827 -1248
rect 247 -1354 271 -1330
rect -351 -1494 -319 -1368
rect -299 -1494 -267 -1368
rect -247 -1432 -215 -1368
rect -195 -1432 -163 -1368
rect -147 -1478 -83 -1414
rect 1250 -1446 1290 -1412
rect 1328 -1451 1352 -1427
rect 1388 -1500 1422 -1464
rect 1429 -1501 1453 -1477
rect 1250 -1551 1290 -1517
rect 1328 -1556 1352 -1532
rect -349 -1720 -317 -1594
rect -297 -1720 -265 -1594
rect -245 -1658 -213 -1594
rect -193 -1658 -161 -1594
rect 1501 -1613 1535 -1577
rect 1542 -1614 1566 -1590
rect -145 -1704 -81 -1640
rect 1250 -1654 1290 -1620
rect 1328 -1659 1352 -1635
rect 1385 -1702 1419 -1666
rect 1426 -1703 1450 -1679
rect 1240 -1743 1280 -1709
rect 1604 -1715 1638 -1679
rect 1645 -1716 1669 -1692
rect 1318 -1748 1342 -1724
rect -349 -1943 -317 -1817
rect -297 -1943 -265 -1817
rect -245 -1881 -213 -1817
rect -193 -1881 -161 -1817
rect -145 -1927 -81 -1863
<< ntransistor >>
rect -217 -362 -215 -342
rect -165 -362 -163 -342
rect -321 -409 -319 -389
rect -269 -409 -267 -389
rect -217 -409 -215 -389
rect -165 -409 -163 -389
rect -117 -392 -115 -372
rect -85 -392 -83 -372
rect 1690 -376 1692 -356
rect 1742 -376 1744 -356
rect 1586 -423 1588 -403
rect 1638 -423 1640 -403
rect 1690 -423 1692 -403
rect 1742 -423 1744 -403
rect 1790 -406 1792 -386
rect 1822 -406 1824 -386
rect 155 -487 157 -483
rect 155 -537 157 -533
rect 186 -537 188 -533
rect 196 -537 198 -533
rect 206 -537 208 -533
rect 216 -537 218 -533
rect -220 -589 -218 -569
rect -168 -589 -166 -569
rect 968 -557 970 -553
rect -324 -636 -322 -616
rect -272 -636 -270 -616
rect -220 -636 -218 -616
rect -168 -636 -166 -616
rect -120 -619 -118 -599
rect -88 -619 -86 -599
rect 156 -608 158 -604
rect 968 -607 970 -603
rect 999 -607 1001 -603
rect 1009 -607 1011 -603
rect 1019 -607 1021 -603
rect 1029 -607 1031 -603
rect 156 -658 158 -654
rect 187 -658 189 -654
rect 197 -658 199 -654
rect 207 -658 209 -654
rect 217 -658 219 -654
rect 1682 -618 1684 -598
rect 1734 -618 1736 -598
rect 720 -673 722 -667
rect 830 -674 832 -668
rect 639 -692 642 -676
rect 652 -692 655 -676
rect 789 -680 791 -674
rect 799 -680 801 -674
rect 978 -681 980 -677
rect 156 -729 158 -725
rect -223 -818 -221 -798
rect -171 -818 -169 -798
rect 1578 -665 1580 -645
rect 1630 -665 1632 -645
rect 1682 -665 1684 -645
rect 1734 -665 1736 -645
rect 1782 -648 1784 -628
rect 1814 -648 1816 -628
rect 978 -731 980 -727
rect 1009 -731 1011 -727
rect 1019 -731 1021 -727
rect 1029 -731 1031 -727
rect 1039 -731 1041 -727
rect 560 -768 562 -758
rect 156 -779 158 -775
rect 187 -779 189 -775
rect 197 -779 199 -775
rect 207 -779 209 -775
rect 217 -779 219 -775
rect 503 -781 505 -771
rect 513 -781 515 -771
rect 521 -781 523 -771
rect 653 -794 655 -788
rect 612 -800 614 -794
rect 622 -800 624 -794
rect -327 -865 -325 -845
rect -275 -865 -273 -845
rect -223 -865 -221 -845
rect -171 -865 -169 -845
rect -123 -848 -121 -828
rect -91 -848 -89 -828
rect 156 -849 158 -845
rect 882 -835 884 -831
rect 576 -864 578 -858
rect 500 -883 503 -867
rect 513 -883 516 -867
rect 156 -899 158 -895
rect 187 -899 189 -895
rect 197 -899 199 -895
rect 207 -899 209 -895
rect 217 -899 219 -895
rect 1683 -854 1685 -834
rect 1735 -854 1737 -834
rect 882 -885 884 -881
rect 913 -885 915 -881
rect 923 -885 925 -881
rect 933 -885 935 -881
rect 943 -885 945 -881
rect 692 -902 694 -896
rect 651 -908 653 -902
rect 661 -908 663 -902
rect 1579 -901 1581 -881
rect 1631 -901 1633 -881
rect 1683 -901 1685 -881
rect 1735 -901 1737 -881
rect 1783 -884 1785 -864
rect 1815 -884 1817 -864
rect -223 -1034 -221 -1014
rect -171 -1034 -169 -1014
rect 935 -1034 937 -1028
rect -327 -1081 -325 -1061
rect -275 -1081 -273 -1061
rect -223 -1081 -221 -1061
rect -171 -1081 -169 -1061
rect -123 -1064 -121 -1044
rect -91 -1064 -89 -1044
rect 858 -1053 861 -1037
rect 871 -1053 874 -1037
rect 254 -1107 256 -1101
rect 177 -1126 180 -1110
rect 190 -1126 193 -1110
rect 1052 -1097 1054 -1091
rect 1011 -1103 1013 -1097
rect 1021 -1103 1023 -1097
rect 1326 -1121 1328 -1117
rect 939 -1141 941 -1135
rect 862 -1160 865 -1144
rect 875 -1160 878 -1144
rect 1683 -1087 1685 -1067
rect 1735 -1087 1737 -1067
rect 1579 -1134 1581 -1114
rect 1631 -1134 1633 -1114
rect 1683 -1134 1685 -1114
rect 1735 -1134 1737 -1114
rect 1783 -1117 1785 -1097
rect 1815 -1117 1817 -1097
rect 1140 -1176 1142 -1170
rect 1326 -1171 1328 -1167
rect 1357 -1171 1359 -1167
rect 1367 -1171 1369 -1167
rect 1377 -1171 1379 -1167
rect 1387 -1171 1389 -1167
rect 1099 -1182 1101 -1176
rect 1109 -1182 1111 -1176
rect 254 -1194 256 -1188
rect -224 -1249 -222 -1229
rect -172 -1249 -170 -1229
rect 178 -1213 181 -1197
rect 191 -1213 194 -1197
rect -328 -1296 -326 -1276
rect -276 -1296 -274 -1276
rect -224 -1296 -222 -1276
rect -172 -1296 -170 -1276
rect -124 -1279 -122 -1259
rect -92 -1279 -90 -1259
rect 939 -1250 941 -1244
rect 862 -1269 865 -1253
rect 875 -1269 878 -1253
rect 1052 -1266 1054 -1260
rect 1011 -1272 1013 -1266
rect 1021 -1272 1023 -1266
rect 257 -1282 259 -1276
rect 180 -1301 183 -1285
rect 193 -1301 196 -1285
rect 1678 -1313 1680 -1293
rect 1730 -1313 1732 -1293
rect 1574 -1360 1576 -1340
rect 1626 -1360 1628 -1340
rect 1678 -1360 1680 -1340
rect 1730 -1360 1732 -1340
rect 1778 -1343 1780 -1323
rect 1810 -1343 1812 -1323
rect 258 -1368 260 -1362
rect 180 -1387 183 -1371
rect 193 -1387 196 -1371
rect -232 -1479 -230 -1459
rect -180 -1479 -178 -1459
rect 1339 -1465 1341 -1459
rect 1262 -1484 1265 -1468
rect 1275 -1484 1278 -1468
rect -336 -1526 -334 -1506
rect -284 -1526 -282 -1506
rect -232 -1526 -230 -1506
rect -180 -1526 -178 -1506
rect -132 -1509 -130 -1489
rect -100 -1509 -98 -1489
rect 1440 -1515 1442 -1509
rect 1399 -1521 1401 -1515
rect 1409 -1521 1411 -1515
rect 1339 -1570 1341 -1564
rect 1262 -1589 1265 -1573
rect 1275 -1589 1278 -1573
rect 1553 -1628 1555 -1622
rect 1512 -1634 1514 -1628
rect 1522 -1634 1524 -1628
rect -230 -1705 -228 -1685
rect -178 -1705 -176 -1685
rect 1339 -1673 1341 -1667
rect 1262 -1692 1265 -1676
rect 1275 -1692 1278 -1676
rect -334 -1752 -332 -1732
rect -282 -1752 -280 -1732
rect -230 -1752 -228 -1732
rect -178 -1752 -176 -1732
rect -130 -1735 -128 -1715
rect -98 -1735 -96 -1715
rect 1437 -1717 1439 -1711
rect 1396 -1723 1398 -1717
rect 1406 -1723 1408 -1717
rect 1656 -1730 1658 -1724
rect 1615 -1736 1617 -1730
rect 1625 -1736 1627 -1730
rect 1329 -1762 1331 -1756
rect 1252 -1781 1255 -1765
rect 1265 -1781 1268 -1765
rect -230 -1928 -228 -1908
rect -178 -1928 -176 -1908
rect -334 -1975 -332 -1955
rect -282 -1975 -280 -1955
rect -230 -1975 -228 -1955
rect -178 -1975 -176 -1955
rect -130 -1958 -128 -1938
rect -98 -1958 -96 -1938
<< ptransistor >>
rect -321 -306 -319 -266
rect -269 -306 -267 -266
rect -217 -306 -215 -266
rect -165 -306 -163 -266
rect -321 -368 -319 -328
rect -269 -368 -267 -328
rect -117 -352 -115 -312
rect -85 -352 -83 -312
rect 1586 -320 1588 -280
rect 1638 -320 1640 -280
rect 1690 -320 1692 -280
rect 1742 -320 1744 -280
rect 1586 -382 1588 -342
rect 1638 -382 1640 -342
rect 1790 -366 1792 -326
rect 1822 -366 1824 -326
rect 155 -469 157 -461
rect 186 -469 188 -461
rect 196 -469 198 -461
rect 206 -469 208 -461
rect 216 -469 218 -461
rect -324 -533 -322 -493
rect -272 -533 -270 -493
rect -220 -533 -218 -493
rect -168 -533 -166 -493
rect 155 -519 157 -511
rect -324 -595 -322 -555
rect -272 -595 -270 -555
rect -120 -579 -118 -539
rect -88 -579 -86 -539
rect 968 -539 970 -531
rect 999 -539 1001 -531
rect 1009 -539 1011 -531
rect 1019 -539 1021 -531
rect 1029 -539 1031 -531
rect 156 -590 158 -582
rect 187 -590 189 -582
rect 197 -590 199 -582
rect 207 -590 209 -582
rect 217 -590 219 -582
rect 156 -640 158 -632
rect 968 -589 970 -581
rect 1578 -562 1580 -522
rect 1630 -562 1632 -522
rect 1682 -562 1684 -522
rect 1734 -562 1736 -522
rect 639 -648 642 -628
rect 652 -648 655 -628
rect 720 -653 722 -641
rect 789 -653 791 -629
rect 799 -653 801 -629
rect 1578 -624 1580 -584
rect 1630 -624 1632 -584
rect 1782 -608 1784 -568
rect 1814 -608 1816 -568
rect 830 -654 832 -642
rect 978 -663 980 -655
rect 1009 -663 1011 -655
rect 1019 -663 1021 -655
rect 1029 -663 1031 -655
rect 1039 -663 1041 -655
rect 156 -711 158 -703
rect 187 -711 189 -703
rect 197 -711 199 -703
rect 207 -711 209 -703
rect 217 -711 219 -703
rect -327 -762 -325 -722
rect -275 -762 -273 -722
rect -223 -762 -221 -722
rect -171 -762 -169 -722
rect 156 -761 158 -753
rect -327 -824 -325 -784
rect -275 -824 -273 -784
rect -123 -808 -121 -768
rect -91 -808 -89 -768
rect 978 -713 980 -705
rect 503 -739 505 -714
rect 513 -739 515 -714
rect 521 -739 523 -714
rect 560 -737 562 -717
rect 612 -773 614 -749
rect 622 -773 624 -749
rect 653 -774 655 -762
rect 1579 -798 1581 -758
rect 1631 -798 1633 -758
rect 1683 -798 1685 -758
rect 1735 -798 1737 -758
rect 156 -831 158 -823
rect 187 -831 189 -823
rect 197 -831 199 -823
rect 207 -831 209 -823
rect 217 -831 219 -823
rect 156 -881 158 -873
rect 882 -817 884 -809
rect 913 -817 915 -809
rect 923 -817 925 -809
rect 933 -817 935 -809
rect 943 -817 945 -809
rect 500 -839 503 -819
rect 513 -839 516 -819
rect 576 -844 578 -832
rect 651 -881 653 -857
rect 661 -881 663 -857
rect 882 -867 884 -859
rect 692 -882 694 -870
rect 1579 -860 1581 -820
rect 1631 -860 1633 -820
rect 1783 -844 1785 -804
rect 1815 -844 1817 -804
rect -327 -978 -325 -938
rect -275 -978 -273 -938
rect -223 -978 -221 -938
rect -171 -978 -169 -938
rect -327 -1040 -325 -1000
rect -275 -1040 -273 -1000
rect -123 -1024 -121 -984
rect -91 -1024 -89 -984
rect 858 -1009 861 -989
rect 871 -1009 874 -989
rect 935 -1014 937 -1002
rect 1579 -1031 1581 -991
rect 1631 -1031 1633 -991
rect 1683 -1031 1685 -991
rect 1735 -1031 1737 -991
rect 177 -1082 180 -1062
rect 190 -1082 193 -1062
rect 254 -1087 256 -1075
rect 1011 -1076 1013 -1052
rect 1021 -1076 1023 -1052
rect 862 -1116 865 -1096
rect 875 -1116 878 -1096
rect 1052 -1077 1054 -1065
rect 1326 -1103 1328 -1095
rect 1357 -1103 1359 -1095
rect 1367 -1103 1369 -1095
rect 1377 -1103 1379 -1095
rect 1387 -1103 1389 -1095
rect 939 -1121 941 -1109
rect -328 -1193 -326 -1153
rect -276 -1193 -274 -1153
rect -224 -1193 -222 -1153
rect -172 -1193 -170 -1153
rect 178 -1169 181 -1149
rect 191 -1169 194 -1149
rect 1099 -1155 1101 -1131
rect 1109 -1155 1111 -1131
rect 254 -1174 256 -1162
rect 1140 -1156 1142 -1144
rect 1326 -1153 1328 -1145
rect 1579 -1093 1581 -1053
rect 1631 -1093 1633 -1053
rect 1783 -1077 1785 -1037
rect 1815 -1077 1817 -1037
rect -328 -1255 -326 -1215
rect -276 -1255 -274 -1215
rect -124 -1239 -122 -1199
rect -92 -1239 -90 -1199
rect 862 -1225 865 -1205
rect 875 -1225 878 -1205
rect 180 -1257 183 -1237
rect 193 -1257 196 -1237
rect 257 -1262 259 -1250
rect 939 -1230 941 -1218
rect 1011 -1245 1013 -1221
rect 1021 -1245 1023 -1221
rect 1052 -1246 1054 -1234
rect 1574 -1257 1576 -1217
rect 1626 -1257 1628 -1217
rect 1678 -1257 1680 -1217
rect 1730 -1257 1732 -1217
rect 1574 -1319 1576 -1279
rect 1626 -1319 1628 -1279
rect 1778 -1303 1780 -1263
rect 1810 -1303 1812 -1263
rect 180 -1343 183 -1323
rect 193 -1343 196 -1323
rect 258 -1348 260 -1336
rect -336 -1423 -334 -1383
rect -284 -1423 -282 -1383
rect -232 -1423 -230 -1383
rect -180 -1423 -178 -1383
rect -336 -1485 -334 -1445
rect -284 -1485 -282 -1445
rect -132 -1469 -130 -1429
rect -100 -1469 -98 -1429
rect 1262 -1440 1265 -1420
rect 1275 -1440 1278 -1420
rect 1339 -1445 1341 -1433
rect 1399 -1494 1401 -1470
rect 1409 -1494 1411 -1470
rect 1440 -1495 1442 -1483
rect 1262 -1545 1265 -1525
rect 1275 -1545 1278 -1525
rect 1339 -1550 1341 -1538
rect 1512 -1607 1514 -1583
rect 1522 -1607 1524 -1583
rect -334 -1649 -332 -1609
rect -282 -1649 -280 -1609
rect -230 -1649 -228 -1609
rect -178 -1649 -176 -1609
rect 1553 -1608 1555 -1596
rect 1262 -1648 1265 -1628
rect 1275 -1648 1278 -1628
rect -334 -1711 -332 -1671
rect -282 -1711 -280 -1671
rect -130 -1695 -128 -1655
rect -98 -1695 -96 -1655
rect 1339 -1653 1341 -1641
rect 1396 -1696 1398 -1672
rect 1406 -1696 1408 -1672
rect 1437 -1697 1439 -1685
rect 1615 -1709 1617 -1685
rect 1625 -1709 1627 -1685
rect 1252 -1737 1255 -1717
rect 1265 -1737 1268 -1717
rect 1656 -1710 1658 -1698
rect 1329 -1742 1331 -1730
rect -334 -1872 -332 -1832
rect -282 -1872 -280 -1832
rect -230 -1872 -228 -1832
rect -178 -1872 -176 -1832
rect -334 -1934 -332 -1894
rect -282 -1934 -280 -1894
rect -130 -1918 -128 -1878
rect -98 -1918 -96 -1878
<< ndiffusion >>
rect -218 -362 -217 -342
rect -215 -362 -214 -342
rect -166 -362 -165 -342
rect -163 -362 -162 -342
rect -322 -409 -321 -389
rect -319 -409 -318 -389
rect -270 -409 -269 -389
rect -267 -409 -266 -389
rect -218 -409 -217 -389
rect -215 -409 -214 -389
rect -166 -409 -165 -389
rect -163 -409 -162 -389
rect -118 -392 -117 -372
rect -115 -392 -114 -372
rect -86 -392 -85 -372
rect -83 -392 -82 -372
rect 1689 -376 1690 -356
rect 1692 -376 1693 -356
rect 1741 -376 1742 -356
rect 1744 -376 1745 -356
rect 1585 -423 1586 -403
rect 1588 -423 1589 -403
rect 1637 -423 1638 -403
rect 1640 -423 1641 -403
rect 1689 -423 1690 -403
rect 1692 -423 1693 -403
rect 1741 -423 1742 -403
rect 1744 -423 1745 -403
rect 1789 -406 1790 -386
rect 1792 -406 1793 -386
rect 1821 -406 1822 -386
rect 1824 -406 1825 -386
rect 154 -487 155 -483
rect 157 -487 158 -483
rect 154 -537 155 -533
rect 157 -537 158 -533
rect 184 -537 186 -533
rect 188 -537 196 -533
rect 198 -537 200 -533
rect 204 -537 206 -533
rect 208 -537 216 -533
rect 218 -537 220 -533
rect -221 -589 -220 -569
rect -218 -589 -217 -569
rect -169 -589 -168 -569
rect -166 -589 -165 -569
rect 967 -557 968 -553
rect 970 -557 971 -553
rect -325 -636 -324 -616
rect -322 -636 -321 -616
rect -273 -636 -272 -616
rect -270 -636 -269 -616
rect -221 -636 -220 -616
rect -218 -636 -217 -616
rect -169 -636 -168 -616
rect -166 -636 -165 -616
rect -121 -619 -120 -599
rect -118 -619 -117 -599
rect -89 -619 -88 -599
rect -86 -619 -85 -599
rect 155 -608 156 -604
rect 158 -608 159 -604
rect 967 -607 968 -603
rect 970 -607 971 -603
rect 997 -607 999 -603
rect 1001 -607 1009 -603
rect 1011 -607 1013 -603
rect 1017 -607 1019 -603
rect 1021 -607 1029 -603
rect 1031 -607 1033 -603
rect 155 -658 156 -654
rect 158 -658 159 -654
rect 185 -658 187 -654
rect 189 -658 197 -654
rect 199 -658 201 -654
rect 205 -658 207 -654
rect 209 -658 217 -654
rect 219 -658 221 -654
rect 1681 -618 1682 -598
rect 1684 -618 1685 -598
rect 1733 -618 1734 -598
rect 1736 -618 1737 -598
rect 719 -673 720 -667
rect 722 -673 723 -667
rect 829 -674 830 -668
rect 832 -674 833 -668
rect 637 -681 639 -676
rect 633 -692 639 -681
rect 642 -692 652 -676
rect 655 -681 657 -676
rect 788 -680 789 -674
rect 791 -680 793 -674
rect 797 -680 799 -674
rect 801 -680 802 -674
rect 655 -692 661 -681
rect 977 -681 978 -677
rect 980 -681 981 -677
rect 155 -729 156 -725
rect 158 -729 159 -725
rect -224 -818 -223 -798
rect -221 -818 -220 -798
rect -172 -818 -171 -798
rect -169 -818 -168 -798
rect 1577 -665 1578 -645
rect 1580 -665 1581 -645
rect 1629 -665 1630 -645
rect 1632 -665 1633 -645
rect 1681 -665 1682 -645
rect 1684 -665 1685 -645
rect 1733 -665 1734 -645
rect 1736 -665 1737 -645
rect 1781 -648 1782 -628
rect 1784 -648 1785 -628
rect 1813 -648 1814 -628
rect 1816 -648 1817 -628
rect 977 -731 978 -727
rect 980 -731 981 -727
rect 1007 -731 1009 -727
rect 1011 -731 1019 -727
rect 1021 -731 1023 -727
rect 1027 -731 1029 -727
rect 1031 -731 1039 -727
rect 1041 -731 1043 -727
rect 554 -762 560 -758
rect 554 -768 555 -762
rect 559 -768 560 -762
rect 562 -762 564 -758
rect 569 -762 570 -758
rect 562 -768 570 -762
rect 155 -779 156 -775
rect 158 -779 159 -775
rect 185 -779 187 -775
rect 189 -779 197 -775
rect 199 -779 201 -775
rect 205 -779 207 -775
rect 209 -779 217 -775
rect 219 -779 221 -775
rect 495 -777 503 -771
rect 495 -781 496 -777
rect 501 -781 503 -777
rect 505 -781 513 -771
rect 515 -781 521 -771
rect 523 -775 527 -771
rect 531 -775 532 -771
rect 523 -781 532 -775
rect 652 -794 653 -788
rect 655 -794 656 -788
rect 611 -800 612 -794
rect 614 -800 616 -794
rect 620 -800 622 -794
rect 624 -800 625 -794
rect -328 -865 -327 -845
rect -325 -865 -324 -845
rect -276 -865 -275 -845
rect -273 -865 -272 -845
rect -224 -865 -223 -845
rect -221 -865 -220 -845
rect -172 -865 -171 -845
rect -169 -865 -168 -845
rect -124 -848 -123 -828
rect -121 -848 -120 -828
rect -92 -848 -91 -828
rect -89 -848 -88 -828
rect 155 -849 156 -845
rect 158 -849 159 -845
rect 881 -835 882 -831
rect 884 -835 885 -831
rect 575 -864 576 -858
rect 578 -864 579 -858
rect 498 -872 500 -867
rect 494 -883 500 -872
rect 503 -883 513 -867
rect 516 -872 518 -867
rect 516 -883 522 -872
rect 155 -899 156 -895
rect 158 -899 159 -895
rect 185 -899 187 -895
rect 189 -899 197 -895
rect 199 -899 201 -895
rect 205 -899 207 -895
rect 209 -899 217 -895
rect 219 -899 221 -895
rect 1682 -854 1683 -834
rect 1685 -854 1686 -834
rect 1734 -854 1735 -834
rect 1737 -854 1738 -834
rect 881 -885 882 -881
rect 884 -885 885 -881
rect 911 -885 913 -881
rect 915 -885 923 -881
rect 925 -885 927 -881
rect 931 -885 933 -881
rect 935 -885 943 -881
rect 945 -885 947 -881
rect 691 -902 692 -896
rect 694 -902 695 -896
rect 650 -908 651 -902
rect 653 -908 655 -902
rect 659 -908 661 -902
rect 663 -908 664 -902
rect 1578 -901 1579 -881
rect 1581 -901 1582 -881
rect 1630 -901 1631 -881
rect 1633 -901 1634 -881
rect 1682 -901 1683 -881
rect 1685 -901 1686 -881
rect 1734 -901 1735 -881
rect 1737 -901 1738 -881
rect 1782 -884 1783 -864
rect 1785 -884 1786 -864
rect 1814 -884 1815 -864
rect 1817 -884 1818 -864
rect -224 -1034 -223 -1014
rect -221 -1034 -220 -1014
rect -172 -1034 -171 -1014
rect -169 -1034 -168 -1014
rect 934 -1034 935 -1028
rect 937 -1034 938 -1028
rect 856 -1042 858 -1037
rect -328 -1081 -327 -1061
rect -325 -1081 -324 -1061
rect -276 -1081 -275 -1061
rect -273 -1081 -272 -1061
rect -224 -1081 -223 -1061
rect -221 -1081 -220 -1061
rect -172 -1081 -171 -1061
rect -169 -1081 -168 -1061
rect -124 -1064 -123 -1044
rect -121 -1064 -120 -1044
rect -92 -1064 -91 -1044
rect -89 -1064 -88 -1044
rect 852 -1053 858 -1042
rect 861 -1053 871 -1037
rect 874 -1042 876 -1037
rect 874 -1053 880 -1042
rect 253 -1107 254 -1101
rect 256 -1107 257 -1101
rect 175 -1115 177 -1110
rect 171 -1126 177 -1115
rect 180 -1126 190 -1110
rect 193 -1115 195 -1110
rect 193 -1126 199 -1115
rect 1051 -1097 1052 -1091
rect 1054 -1097 1055 -1091
rect 1010 -1103 1011 -1097
rect 1013 -1103 1015 -1097
rect 1019 -1103 1021 -1097
rect 1023 -1103 1024 -1097
rect 1325 -1121 1326 -1117
rect 1328 -1121 1329 -1117
rect 938 -1141 939 -1135
rect 941 -1141 942 -1135
rect 860 -1149 862 -1144
rect 856 -1160 862 -1149
rect 865 -1160 875 -1144
rect 878 -1149 880 -1144
rect 878 -1160 884 -1149
rect 1682 -1087 1683 -1067
rect 1685 -1087 1686 -1067
rect 1734 -1087 1735 -1067
rect 1737 -1087 1738 -1067
rect 1578 -1134 1579 -1114
rect 1581 -1134 1582 -1114
rect 1630 -1134 1631 -1114
rect 1633 -1134 1634 -1114
rect 1682 -1134 1683 -1114
rect 1685 -1134 1686 -1114
rect 1734 -1134 1735 -1114
rect 1737 -1134 1738 -1114
rect 1782 -1117 1783 -1097
rect 1785 -1117 1786 -1097
rect 1814 -1117 1815 -1097
rect 1817 -1117 1818 -1097
rect 1139 -1176 1140 -1170
rect 1142 -1176 1143 -1170
rect 1325 -1171 1326 -1167
rect 1328 -1171 1329 -1167
rect 1355 -1171 1357 -1167
rect 1359 -1171 1367 -1167
rect 1369 -1171 1371 -1167
rect 1375 -1171 1377 -1167
rect 1379 -1171 1387 -1167
rect 1389 -1171 1391 -1167
rect 1098 -1182 1099 -1176
rect 1101 -1182 1103 -1176
rect 1107 -1182 1109 -1176
rect 1111 -1182 1112 -1176
rect 253 -1194 254 -1188
rect 256 -1194 257 -1188
rect -225 -1249 -224 -1229
rect -222 -1249 -221 -1229
rect -173 -1249 -172 -1229
rect -170 -1249 -169 -1229
rect 176 -1202 178 -1197
rect 172 -1213 178 -1202
rect 181 -1213 191 -1197
rect 194 -1202 196 -1197
rect 194 -1213 200 -1202
rect -329 -1296 -328 -1276
rect -326 -1296 -325 -1276
rect -277 -1296 -276 -1276
rect -274 -1296 -273 -1276
rect -225 -1296 -224 -1276
rect -222 -1296 -221 -1276
rect -173 -1296 -172 -1276
rect -170 -1296 -169 -1276
rect -125 -1279 -124 -1259
rect -122 -1279 -121 -1259
rect -93 -1279 -92 -1259
rect -90 -1279 -89 -1259
rect 938 -1250 939 -1244
rect 941 -1250 942 -1244
rect 860 -1258 862 -1253
rect 856 -1269 862 -1258
rect 865 -1269 875 -1253
rect 878 -1258 880 -1253
rect 878 -1269 884 -1258
rect 1051 -1266 1052 -1260
rect 1054 -1266 1055 -1260
rect 1010 -1272 1011 -1266
rect 1013 -1272 1015 -1266
rect 1019 -1272 1021 -1266
rect 1023 -1272 1024 -1266
rect 256 -1282 257 -1276
rect 259 -1282 260 -1276
rect 178 -1290 180 -1285
rect 174 -1301 180 -1290
rect 183 -1301 193 -1285
rect 196 -1290 198 -1285
rect 196 -1301 202 -1290
rect 1677 -1313 1678 -1293
rect 1680 -1313 1681 -1293
rect 1729 -1313 1730 -1293
rect 1732 -1313 1733 -1293
rect 1573 -1360 1574 -1340
rect 1576 -1360 1577 -1340
rect 1625 -1360 1626 -1340
rect 1628 -1360 1629 -1340
rect 1677 -1360 1678 -1340
rect 1680 -1360 1681 -1340
rect 1729 -1360 1730 -1340
rect 1732 -1360 1733 -1340
rect 1777 -1343 1778 -1323
rect 1780 -1343 1781 -1323
rect 1809 -1343 1810 -1323
rect 1812 -1343 1813 -1323
rect 257 -1368 258 -1362
rect 260 -1368 261 -1362
rect 178 -1376 180 -1371
rect 174 -1387 180 -1376
rect 183 -1387 193 -1371
rect 196 -1376 198 -1371
rect 196 -1387 202 -1376
rect -233 -1479 -232 -1459
rect -230 -1479 -229 -1459
rect -181 -1479 -180 -1459
rect -178 -1479 -177 -1459
rect 1338 -1465 1339 -1459
rect 1341 -1465 1342 -1459
rect 1260 -1473 1262 -1468
rect 1256 -1484 1262 -1473
rect 1265 -1484 1275 -1468
rect 1278 -1473 1280 -1468
rect 1278 -1484 1284 -1473
rect -337 -1526 -336 -1506
rect -334 -1526 -333 -1506
rect -285 -1526 -284 -1506
rect -282 -1526 -281 -1506
rect -233 -1526 -232 -1506
rect -230 -1526 -229 -1506
rect -181 -1526 -180 -1506
rect -178 -1526 -177 -1506
rect -133 -1509 -132 -1489
rect -130 -1509 -129 -1489
rect -101 -1509 -100 -1489
rect -98 -1509 -97 -1489
rect 1439 -1515 1440 -1509
rect 1442 -1515 1443 -1509
rect 1398 -1521 1399 -1515
rect 1401 -1521 1403 -1515
rect 1407 -1521 1409 -1515
rect 1411 -1521 1412 -1515
rect 1338 -1570 1339 -1564
rect 1341 -1570 1342 -1564
rect 1260 -1578 1262 -1573
rect 1256 -1589 1262 -1578
rect 1265 -1589 1275 -1573
rect 1278 -1578 1280 -1573
rect 1278 -1589 1284 -1578
rect 1552 -1628 1553 -1622
rect 1555 -1628 1556 -1622
rect 1511 -1634 1512 -1628
rect 1514 -1634 1516 -1628
rect 1520 -1634 1522 -1628
rect 1524 -1634 1525 -1628
rect -231 -1705 -230 -1685
rect -228 -1705 -227 -1685
rect -179 -1705 -178 -1685
rect -176 -1705 -175 -1685
rect 1338 -1673 1339 -1667
rect 1341 -1673 1342 -1667
rect 1260 -1681 1262 -1676
rect 1256 -1692 1262 -1681
rect 1265 -1692 1275 -1676
rect 1278 -1681 1280 -1676
rect 1278 -1692 1284 -1681
rect -335 -1752 -334 -1732
rect -332 -1752 -331 -1732
rect -283 -1752 -282 -1732
rect -280 -1752 -279 -1732
rect -231 -1752 -230 -1732
rect -228 -1752 -227 -1732
rect -179 -1752 -178 -1732
rect -176 -1752 -175 -1732
rect -131 -1735 -130 -1715
rect -128 -1735 -127 -1715
rect -99 -1735 -98 -1715
rect -96 -1735 -95 -1715
rect 1436 -1717 1437 -1711
rect 1439 -1717 1440 -1711
rect 1395 -1723 1396 -1717
rect 1398 -1723 1400 -1717
rect 1404 -1723 1406 -1717
rect 1408 -1723 1409 -1717
rect 1655 -1730 1656 -1724
rect 1658 -1730 1659 -1724
rect 1614 -1736 1615 -1730
rect 1617 -1736 1619 -1730
rect 1623 -1736 1625 -1730
rect 1627 -1736 1628 -1730
rect 1328 -1762 1329 -1756
rect 1331 -1762 1332 -1756
rect 1250 -1770 1252 -1765
rect 1246 -1781 1252 -1770
rect 1255 -1781 1265 -1765
rect 1268 -1770 1270 -1765
rect 1268 -1781 1274 -1770
rect -231 -1928 -230 -1908
rect -228 -1928 -227 -1908
rect -179 -1928 -178 -1908
rect -176 -1928 -175 -1908
rect -335 -1975 -334 -1955
rect -332 -1975 -331 -1955
rect -283 -1975 -282 -1955
rect -280 -1975 -279 -1955
rect -231 -1975 -230 -1955
rect -228 -1975 -227 -1955
rect -179 -1975 -178 -1955
rect -176 -1975 -175 -1955
rect -131 -1958 -130 -1938
rect -128 -1958 -127 -1938
rect -99 -1958 -98 -1938
rect -96 -1958 -95 -1938
<< pdiffusion >>
rect -322 -306 -321 -266
rect -319 -306 -318 -266
rect -270 -306 -269 -266
rect -267 -306 -266 -266
rect -218 -306 -217 -266
rect -215 -306 -214 -266
rect -166 -306 -165 -266
rect -163 -306 -162 -266
rect -322 -368 -321 -328
rect -319 -368 -318 -328
rect -270 -368 -269 -328
rect -267 -368 -266 -328
rect -118 -352 -117 -312
rect -115 -352 -114 -312
rect -86 -352 -85 -312
rect -83 -352 -82 -312
rect 1585 -320 1586 -280
rect 1588 -320 1589 -280
rect 1637 -320 1638 -280
rect 1640 -320 1641 -280
rect 1689 -320 1690 -280
rect 1692 -320 1693 -280
rect 1741 -320 1742 -280
rect 1744 -320 1745 -280
rect 1585 -382 1586 -342
rect 1588 -382 1589 -342
rect 1637 -382 1638 -342
rect 1640 -382 1641 -342
rect 1789 -366 1790 -326
rect 1792 -366 1793 -326
rect 1821 -366 1822 -326
rect 1824 -366 1825 -326
rect 154 -469 155 -461
rect 157 -469 158 -461
rect 184 -469 186 -461
rect 188 -469 196 -461
rect 198 -469 200 -461
rect 204 -469 206 -461
rect 208 -469 216 -461
rect 218 -469 220 -461
rect -325 -533 -324 -493
rect -322 -533 -321 -493
rect -273 -533 -272 -493
rect -270 -533 -269 -493
rect -221 -533 -220 -493
rect -218 -533 -217 -493
rect -169 -533 -168 -493
rect -166 -533 -165 -493
rect 154 -519 155 -511
rect 157 -519 158 -511
rect -325 -595 -324 -555
rect -322 -595 -321 -555
rect -273 -595 -272 -555
rect -270 -595 -269 -555
rect -121 -579 -120 -539
rect -118 -579 -117 -539
rect -89 -579 -88 -539
rect -86 -579 -85 -539
rect 967 -539 968 -531
rect 970 -539 971 -531
rect 997 -539 999 -531
rect 1001 -539 1009 -531
rect 1011 -539 1013 -531
rect 1017 -539 1019 -531
rect 1021 -539 1029 -531
rect 1031 -539 1033 -531
rect 155 -590 156 -582
rect 158 -590 159 -582
rect 185 -590 187 -582
rect 189 -590 197 -582
rect 199 -590 201 -582
rect 205 -590 207 -582
rect 209 -590 217 -582
rect 219 -590 221 -582
rect 155 -640 156 -632
rect 158 -640 159 -632
rect 967 -589 968 -581
rect 970 -589 971 -581
rect 1577 -562 1578 -522
rect 1580 -562 1581 -522
rect 1629 -562 1630 -522
rect 1632 -562 1633 -522
rect 1681 -562 1682 -522
rect 1684 -562 1685 -522
rect 1733 -562 1734 -522
rect 1736 -562 1737 -522
rect 637 -633 639 -628
rect 633 -648 639 -633
rect 642 -633 645 -628
rect 649 -633 652 -628
rect 642 -648 652 -633
rect 655 -633 657 -628
rect 655 -648 661 -633
rect 719 -653 720 -641
rect 722 -653 723 -641
rect 788 -653 789 -629
rect 791 -653 799 -629
rect 801 -653 802 -629
rect 1577 -624 1578 -584
rect 1580 -624 1581 -584
rect 1629 -624 1630 -584
rect 1632 -624 1633 -584
rect 1781 -608 1782 -568
rect 1784 -608 1785 -568
rect 1813 -608 1814 -568
rect 1816 -608 1817 -568
rect 829 -654 830 -642
rect 832 -654 833 -642
rect 977 -663 978 -655
rect 980 -663 981 -655
rect 1007 -663 1009 -655
rect 1011 -663 1019 -655
rect 1021 -663 1023 -655
rect 1027 -663 1029 -655
rect 1031 -663 1039 -655
rect 1041 -663 1043 -655
rect 155 -711 156 -703
rect 158 -711 159 -703
rect 185 -711 187 -703
rect 189 -711 197 -703
rect 199 -711 201 -703
rect 205 -711 207 -703
rect 209 -711 217 -703
rect 219 -711 221 -703
rect -328 -762 -327 -722
rect -325 -762 -324 -722
rect -276 -762 -275 -722
rect -273 -762 -272 -722
rect -224 -762 -223 -722
rect -221 -762 -220 -722
rect -172 -762 -171 -722
rect -169 -762 -168 -722
rect 155 -761 156 -753
rect 158 -761 159 -753
rect -328 -824 -327 -784
rect -325 -824 -324 -784
rect -276 -824 -275 -784
rect -273 -824 -272 -784
rect -124 -808 -123 -768
rect -121 -808 -120 -768
rect -92 -808 -91 -768
rect -89 -808 -88 -768
rect 977 -713 978 -705
rect 980 -713 981 -705
rect 495 -718 496 -714
rect 500 -718 503 -714
rect 495 -739 503 -718
rect 505 -735 513 -714
rect 505 -739 507 -735
rect 511 -739 513 -735
rect 515 -718 516 -714
rect 520 -718 521 -714
rect 515 -739 521 -718
rect 523 -734 532 -714
rect 523 -739 527 -734
rect 531 -739 532 -734
rect 559 -724 560 -717
rect 554 -737 560 -724
rect 562 -732 570 -717
rect 562 -737 564 -732
rect 569 -737 570 -732
rect 611 -773 612 -749
rect 614 -773 622 -749
rect 624 -773 625 -749
rect 652 -774 653 -762
rect 655 -774 656 -762
rect 1578 -798 1579 -758
rect 1581 -798 1582 -758
rect 1630 -798 1631 -758
rect 1633 -798 1634 -758
rect 1682 -798 1683 -758
rect 1685 -798 1686 -758
rect 1734 -798 1735 -758
rect 1737 -798 1738 -758
rect 155 -831 156 -823
rect 158 -831 159 -823
rect 185 -831 187 -823
rect 189 -831 197 -823
rect 199 -831 201 -823
rect 205 -831 207 -823
rect 209 -831 217 -823
rect 219 -831 221 -823
rect 155 -881 156 -873
rect 158 -881 159 -873
rect 881 -817 882 -809
rect 884 -817 885 -809
rect 911 -817 913 -809
rect 915 -817 923 -809
rect 925 -817 927 -809
rect 931 -817 933 -809
rect 935 -817 943 -809
rect 945 -817 947 -809
rect 498 -824 500 -819
rect 494 -839 500 -824
rect 503 -824 506 -819
rect 510 -824 513 -819
rect 503 -839 513 -824
rect 516 -824 518 -819
rect 516 -839 522 -824
rect 575 -844 576 -832
rect 578 -844 579 -832
rect 650 -881 651 -857
rect 653 -881 661 -857
rect 663 -881 664 -857
rect 881 -867 882 -859
rect 884 -867 885 -859
rect 691 -882 692 -870
rect 694 -882 695 -870
rect 1578 -860 1579 -820
rect 1581 -860 1582 -820
rect 1630 -860 1631 -820
rect 1633 -860 1634 -820
rect 1782 -844 1783 -804
rect 1785 -844 1786 -804
rect 1814 -844 1815 -804
rect 1817 -844 1818 -804
rect -328 -978 -327 -938
rect -325 -978 -324 -938
rect -276 -978 -275 -938
rect -273 -978 -272 -938
rect -224 -978 -223 -938
rect -221 -978 -220 -938
rect -172 -978 -171 -938
rect -169 -978 -168 -938
rect -328 -1040 -327 -1000
rect -325 -1040 -324 -1000
rect -276 -1040 -275 -1000
rect -273 -1040 -272 -1000
rect -124 -1024 -123 -984
rect -121 -1024 -120 -984
rect -92 -1024 -91 -984
rect -89 -1024 -88 -984
rect 856 -994 858 -989
rect 852 -1009 858 -994
rect 861 -994 864 -989
rect 868 -994 871 -989
rect 861 -1009 871 -994
rect 874 -994 876 -989
rect 874 -1009 880 -994
rect 934 -1014 935 -1002
rect 937 -1014 938 -1002
rect 1578 -1031 1579 -991
rect 1581 -1031 1582 -991
rect 1630 -1031 1631 -991
rect 1633 -1031 1634 -991
rect 1682 -1031 1683 -991
rect 1685 -1031 1686 -991
rect 1734 -1031 1735 -991
rect 1737 -1031 1738 -991
rect 175 -1067 177 -1062
rect 171 -1082 177 -1067
rect 180 -1067 183 -1062
rect 187 -1067 190 -1062
rect 180 -1082 190 -1067
rect 193 -1067 195 -1062
rect 193 -1082 199 -1067
rect 253 -1087 254 -1075
rect 256 -1087 257 -1075
rect 1010 -1076 1011 -1052
rect 1013 -1076 1021 -1052
rect 1023 -1076 1024 -1052
rect 860 -1101 862 -1096
rect 856 -1116 862 -1101
rect 865 -1101 868 -1096
rect 872 -1101 875 -1096
rect 865 -1116 875 -1101
rect 878 -1101 880 -1096
rect 1051 -1077 1052 -1065
rect 1054 -1077 1055 -1065
rect 878 -1116 884 -1101
rect 1325 -1103 1326 -1095
rect 1328 -1103 1329 -1095
rect 1355 -1103 1357 -1095
rect 1359 -1103 1367 -1095
rect 1369 -1103 1371 -1095
rect 1375 -1103 1377 -1095
rect 1379 -1103 1387 -1095
rect 1389 -1103 1391 -1095
rect 938 -1121 939 -1109
rect 941 -1121 942 -1109
rect -329 -1193 -328 -1153
rect -326 -1193 -325 -1153
rect -277 -1193 -276 -1153
rect -274 -1193 -273 -1153
rect -225 -1193 -224 -1153
rect -222 -1193 -221 -1153
rect -173 -1193 -172 -1153
rect -170 -1193 -169 -1153
rect 176 -1154 178 -1149
rect 172 -1169 178 -1154
rect 181 -1154 184 -1149
rect 188 -1154 191 -1149
rect 181 -1169 191 -1154
rect 194 -1154 196 -1149
rect 194 -1169 200 -1154
rect 1098 -1155 1099 -1131
rect 1101 -1155 1109 -1131
rect 1111 -1155 1112 -1131
rect 253 -1174 254 -1162
rect 256 -1174 257 -1162
rect 1139 -1156 1140 -1144
rect 1142 -1156 1143 -1144
rect 1325 -1153 1326 -1145
rect 1328 -1153 1329 -1145
rect 1578 -1093 1579 -1053
rect 1581 -1093 1582 -1053
rect 1630 -1093 1631 -1053
rect 1633 -1093 1634 -1053
rect 1782 -1077 1783 -1037
rect 1785 -1077 1786 -1037
rect 1814 -1077 1815 -1037
rect 1817 -1077 1818 -1037
rect -329 -1255 -328 -1215
rect -326 -1255 -325 -1215
rect -277 -1255 -276 -1215
rect -274 -1255 -273 -1215
rect -125 -1239 -124 -1199
rect -122 -1239 -121 -1199
rect -93 -1239 -92 -1199
rect -90 -1239 -89 -1199
rect 860 -1210 862 -1205
rect 856 -1225 862 -1210
rect 865 -1210 868 -1205
rect 872 -1210 875 -1205
rect 865 -1225 875 -1210
rect 878 -1210 880 -1205
rect 878 -1225 884 -1210
rect 178 -1242 180 -1237
rect 174 -1257 180 -1242
rect 183 -1242 186 -1237
rect 190 -1242 193 -1237
rect 183 -1257 193 -1242
rect 196 -1242 198 -1237
rect 196 -1257 202 -1242
rect 256 -1262 257 -1250
rect 259 -1262 260 -1250
rect 938 -1230 939 -1218
rect 941 -1230 942 -1218
rect 1010 -1245 1011 -1221
rect 1013 -1245 1021 -1221
rect 1023 -1245 1024 -1221
rect 1051 -1246 1052 -1234
rect 1054 -1246 1055 -1234
rect 1573 -1257 1574 -1217
rect 1576 -1257 1577 -1217
rect 1625 -1257 1626 -1217
rect 1628 -1257 1629 -1217
rect 1677 -1257 1678 -1217
rect 1680 -1257 1681 -1217
rect 1729 -1257 1730 -1217
rect 1732 -1257 1733 -1217
rect 1573 -1319 1574 -1279
rect 1576 -1319 1577 -1279
rect 1625 -1319 1626 -1279
rect 1628 -1319 1629 -1279
rect 1777 -1303 1778 -1263
rect 1780 -1303 1781 -1263
rect 1809 -1303 1810 -1263
rect 1812 -1303 1813 -1263
rect 178 -1328 180 -1323
rect 174 -1343 180 -1328
rect 183 -1328 186 -1323
rect 190 -1328 193 -1323
rect 183 -1343 193 -1328
rect 196 -1328 198 -1323
rect 196 -1343 202 -1328
rect 257 -1348 258 -1336
rect 260 -1348 261 -1336
rect -337 -1423 -336 -1383
rect -334 -1423 -333 -1383
rect -285 -1423 -284 -1383
rect -282 -1423 -281 -1383
rect -233 -1423 -232 -1383
rect -230 -1423 -229 -1383
rect -181 -1423 -180 -1383
rect -178 -1423 -177 -1383
rect 1260 -1425 1262 -1420
rect -337 -1485 -336 -1445
rect -334 -1485 -333 -1445
rect -285 -1485 -284 -1445
rect -282 -1485 -281 -1445
rect -133 -1469 -132 -1429
rect -130 -1469 -129 -1429
rect -101 -1469 -100 -1429
rect -98 -1469 -97 -1429
rect 1256 -1440 1262 -1425
rect 1265 -1425 1268 -1420
rect 1272 -1425 1275 -1420
rect 1265 -1440 1275 -1425
rect 1278 -1425 1280 -1420
rect 1278 -1440 1284 -1425
rect 1338 -1445 1339 -1433
rect 1341 -1445 1342 -1433
rect 1398 -1494 1399 -1470
rect 1401 -1494 1409 -1470
rect 1411 -1494 1412 -1470
rect 1439 -1495 1440 -1483
rect 1442 -1495 1443 -1483
rect 1260 -1530 1262 -1525
rect 1256 -1545 1262 -1530
rect 1265 -1530 1268 -1525
rect 1272 -1530 1275 -1525
rect 1265 -1545 1275 -1530
rect 1278 -1530 1280 -1525
rect 1278 -1545 1284 -1530
rect 1338 -1550 1339 -1538
rect 1341 -1550 1342 -1538
rect 1511 -1607 1512 -1583
rect 1514 -1607 1522 -1583
rect 1524 -1607 1525 -1583
rect -335 -1649 -334 -1609
rect -332 -1649 -331 -1609
rect -283 -1649 -282 -1609
rect -280 -1649 -279 -1609
rect -231 -1649 -230 -1609
rect -228 -1649 -227 -1609
rect -179 -1649 -178 -1609
rect -176 -1649 -175 -1609
rect 1552 -1608 1553 -1596
rect 1555 -1608 1556 -1596
rect 1260 -1633 1262 -1628
rect 1256 -1648 1262 -1633
rect 1265 -1633 1268 -1628
rect 1272 -1633 1275 -1628
rect 1265 -1648 1275 -1633
rect 1278 -1633 1280 -1628
rect 1278 -1648 1284 -1633
rect -335 -1711 -334 -1671
rect -332 -1711 -331 -1671
rect -283 -1711 -282 -1671
rect -280 -1711 -279 -1671
rect -131 -1695 -130 -1655
rect -128 -1695 -127 -1655
rect -99 -1695 -98 -1655
rect -96 -1695 -95 -1655
rect 1338 -1653 1339 -1641
rect 1341 -1653 1342 -1641
rect 1395 -1696 1396 -1672
rect 1398 -1696 1406 -1672
rect 1408 -1696 1409 -1672
rect 1436 -1697 1437 -1685
rect 1439 -1697 1440 -1685
rect 1614 -1709 1615 -1685
rect 1617 -1709 1625 -1685
rect 1627 -1709 1628 -1685
rect 1250 -1722 1252 -1717
rect 1246 -1737 1252 -1722
rect 1255 -1722 1258 -1717
rect 1262 -1722 1265 -1717
rect 1255 -1737 1265 -1722
rect 1268 -1722 1270 -1717
rect 1268 -1737 1274 -1722
rect 1655 -1710 1656 -1698
rect 1658 -1710 1659 -1698
rect 1328 -1742 1329 -1730
rect 1331 -1742 1332 -1730
rect -335 -1872 -334 -1832
rect -332 -1872 -331 -1832
rect -283 -1872 -282 -1832
rect -280 -1872 -279 -1832
rect -231 -1872 -230 -1832
rect -228 -1872 -227 -1832
rect -179 -1872 -178 -1832
rect -176 -1872 -175 -1832
rect -335 -1934 -334 -1894
rect -332 -1934 -331 -1894
rect -283 -1934 -282 -1894
rect -280 -1934 -279 -1894
rect -131 -1918 -130 -1878
rect -128 -1918 -127 -1878
rect -99 -1918 -98 -1878
rect -96 -1918 -95 -1878
<< ndcontact >>
rect -222 -362 -218 -342
rect -214 -362 -210 -342
rect -170 -362 -166 -342
rect -162 -362 -158 -342
rect -326 -409 -322 -389
rect -318 -409 -314 -389
rect -274 -409 -270 -389
rect -266 -409 -262 -389
rect -222 -409 -218 -389
rect -214 -409 -210 -389
rect -170 -409 -166 -389
rect -162 -409 -158 -389
rect -122 -392 -118 -372
rect -114 -392 -110 -372
rect -90 -392 -86 -372
rect -82 -392 -78 -372
rect 1685 -376 1689 -356
rect 1693 -376 1697 -356
rect 1737 -376 1741 -356
rect 1745 -376 1749 -356
rect 1581 -423 1585 -403
rect 1589 -423 1593 -403
rect 1633 -423 1637 -403
rect 1641 -423 1645 -403
rect 1685 -423 1689 -403
rect 1693 -423 1697 -403
rect 1737 -423 1741 -403
rect 1745 -423 1749 -403
rect 1785 -406 1789 -386
rect 1793 -406 1797 -386
rect 1817 -406 1821 -386
rect 1825 -406 1829 -386
rect 150 -487 154 -483
rect 158 -487 162 -483
rect 150 -537 154 -533
rect 158 -537 162 -533
rect 180 -537 184 -533
rect 200 -537 204 -533
rect 220 -537 224 -533
rect -225 -589 -221 -569
rect -217 -589 -213 -569
rect -173 -589 -169 -569
rect -165 -589 -161 -569
rect 963 -557 967 -553
rect 971 -557 975 -553
rect -329 -636 -325 -616
rect -321 -636 -317 -616
rect -277 -636 -273 -616
rect -269 -636 -265 -616
rect -225 -636 -221 -616
rect -217 -636 -213 -616
rect -173 -636 -169 -616
rect -165 -636 -161 -616
rect -125 -619 -121 -599
rect -117 -619 -113 -599
rect -93 -619 -89 -599
rect -85 -619 -81 -599
rect 151 -608 155 -604
rect 159 -608 163 -604
rect 963 -607 967 -603
rect 971 -607 975 -603
rect 993 -607 997 -603
rect 1013 -607 1017 -603
rect 1033 -607 1037 -603
rect 151 -658 155 -654
rect 159 -658 163 -654
rect 181 -658 185 -654
rect 201 -658 205 -654
rect 221 -658 225 -654
rect 1677 -618 1681 -598
rect 1685 -618 1689 -598
rect 1729 -618 1733 -598
rect 1737 -618 1741 -598
rect 715 -673 719 -667
rect 723 -673 727 -667
rect 825 -674 829 -668
rect 833 -674 837 -668
rect 633 -681 637 -676
rect 657 -681 661 -676
rect 784 -680 788 -674
rect 793 -680 797 -674
rect 802 -680 806 -674
rect 973 -681 977 -677
rect 981 -681 985 -677
rect 151 -729 155 -725
rect 159 -729 163 -725
rect -228 -818 -224 -798
rect -220 -818 -216 -798
rect -176 -818 -172 -798
rect -168 -818 -164 -798
rect 1573 -665 1577 -645
rect 1581 -665 1585 -645
rect 1625 -665 1629 -645
rect 1633 -665 1637 -645
rect 1677 -665 1681 -645
rect 1685 -665 1689 -645
rect 1729 -665 1733 -645
rect 1737 -665 1741 -645
rect 1777 -648 1781 -628
rect 1785 -648 1789 -628
rect 1809 -648 1813 -628
rect 1817 -648 1821 -628
rect 973 -731 977 -727
rect 981 -731 985 -727
rect 1003 -731 1007 -727
rect 1023 -731 1027 -727
rect 1043 -731 1047 -727
rect 555 -768 559 -762
rect 564 -762 569 -758
rect 151 -779 155 -775
rect 159 -779 163 -775
rect 181 -779 185 -775
rect 201 -779 205 -775
rect 221 -779 225 -775
rect 496 -781 501 -777
rect 527 -775 531 -771
rect 648 -794 652 -788
rect 656 -794 660 -788
rect 607 -800 611 -794
rect 616 -800 620 -794
rect 625 -800 629 -794
rect -332 -865 -328 -845
rect -324 -865 -320 -845
rect -280 -865 -276 -845
rect -272 -865 -268 -845
rect -228 -865 -224 -845
rect -220 -865 -216 -845
rect -176 -865 -172 -845
rect -168 -865 -164 -845
rect -128 -848 -124 -828
rect -120 -848 -116 -828
rect -96 -848 -92 -828
rect -88 -848 -84 -828
rect 151 -849 155 -845
rect 159 -849 163 -845
rect 877 -835 881 -831
rect 885 -835 889 -831
rect 571 -864 575 -858
rect 579 -864 583 -858
rect 494 -872 498 -867
rect 518 -872 522 -867
rect 151 -899 155 -895
rect 159 -899 163 -895
rect 181 -899 185 -895
rect 201 -899 205 -895
rect 221 -899 225 -895
rect 1678 -854 1682 -834
rect 1686 -854 1690 -834
rect 1730 -854 1734 -834
rect 1738 -854 1742 -834
rect 877 -885 881 -881
rect 885 -885 889 -881
rect 907 -885 911 -881
rect 927 -885 931 -881
rect 947 -885 951 -881
rect 687 -902 691 -896
rect 695 -902 699 -896
rect 646 -908 650 -902
rect 655 -908 659 -902
rect 664 -908 668 -902
rect 1574 -901 1578 -881
rect 1582 -901 1586 -881
rect 1626 -901 1630 -881
rect 1634 -901 1638 -881
rect 1678 -901 1682 -881
rect 1686 -901 1690 -881
rect 1730 -901 1734 -881
rect 1738 -901 1742 -881
rect 1778 -884 1782 -864
rect 1786 -884 1790 -864
rect 1810 -884 1814 -864
rect 1818 -884 1822 -864
rect -228 -1034 -224 -1014
rect -220 -1034 -216 -1014
rect -176 -1034 -172 -1014
rect -168 -1034 -164 -1014
rect 930 -1034 934 -1028
rect 938 -1034 942 -1028
rect 852 -1042 856 -1037
rect -332 -1081 -328 -1061
rect -324 -1081 -320 -1061
rect -280 -1081 -276 -1061
rect -272 -1081 -268 -1061
rect -228 -1081 -224 -1061
rect -220 -1081 -216 -1061
rect -176 -1081 -172 -1061
rect -168 -1081 -164 -1061
rect -128 -1064 -124 -1044
rect -120 -1064 -116 -1044
rect -96 -1064 -92 -1044
rect -88 -1064 -84 -1044
rect 876 -1042 880 -1037
rect 249 -1107 253 -1101
rect 257 -1107 261 -1101
rect 171 -1115 175 -1110
rect 195 -1115 199 -1110
rect 1047 -1097 1051 -1091
rect 1055 -1097 1059 -1091
rect 1006 -1103 1010 -1097
rect 1015 -1103 1019 -1097
rect 1024 -1103 1028 -1097
rect 1321 -1121 1325 -1117
rect 1329 -1121 1333 -1117
rect 934 -1141 938 -1135
rect 942 -1141 946 -1135
rect 856 -1149 860 -1144
rect 880 -1149 884 -1144
rect 1678 -1087 1682 -1067
rect 1686 -1087 1690 -1067
rect 1730 -1087 1734 -1067
rect 1738 -1087 1742 -1067
rect 1574 -1134 1578 -1114
rect 1582 -1134 1586 -1114
rect 1626 -1134 1630 -1114
rect 1634 -1134 1638 -1114
rect 1678 -1134 1682 -1114
rect 1686 -1134 1690 -1114
rect 1730 -1134 1734 -1114
rect 1738 -1134 1742 -1114
rect 1778 -1117 1782 -1097
rect 1786 -1117 1790 -1097
rect 1810 -1117 1814 -1097
rect 1818 -1117 1822 -1097
rect 1135 -1176 1139 -1170
rect 1143 -1176 1147 -1170
rect 1321 -1171 1325 -1167
rect 1329 -1171 1333 -1167
rect 1351 -1171 1355 -1167
rect 1371 -1171 1375 -1167
rect 1391 -1171 1395 -1167
rect 1094 -1182 1098 -1176
rect 1103 -1182 1107 -1176
rect 1112 -1182 1116 -1176
rect 249 -1194 253 -1188
rect 257 -1194 261 -1188
rect -229 -1249 -225 -1229
rect -221 -1249 -217 -1229
rect -177 -1249 -173 -1229
rect -169 -1249 -165 -1229
rect 172 -1202 176 -1197
rect 196 -1202 200 -1197
rect -333 -1296 -329 -1276
rect -325 -1296 -321 -1276
rect -281 -1296 -277 -1276
rect -273 -1296 -269 -1276
rect -229 -1296 -225 -1276
rect -221 -1296 -217 -1276
rect -177 -1296 -173 -1276
rect -169 -1296 -165 -1276
rect -129 -1279 -125 -1259
rect -121 -1279 -117 -1259
rect -97 -1279 -93 -1259
rect -89 -1279 -85 -1259
rect 934 -1250 938 -1244
rect 942 -1250 946 -1244
rect 856 -1258 860 -1253
rect 880 -1258 884 -1253
rect 1047 -1266 1051 -1260
rect 1055 -1266 1059 -1260
rect 1006 -1272 1010 -1266
rect 1015 -1272 1019 -1266
rect 1024 -1272 1028 -1266
rect 252 -1282 256 -1276
rect 260 -1282 264 -1276
rect 174 -1290 178 -1285
rect 198 -1290 202 -1285
rect 1673 -1313 1677 -1293
rect 1681 -1313 1685 -1293
rect 1725 -1313 1729 -1293
rect 1733 -1313 1737 -1293
rect 1569 -1360 1573 -1340
rect 1577 -1360 1581 -1340
rect 1621 -1360 1625 -1340
rect 1629 -1360 1633 -1340
rect 1673 -1360 1677 -1340
rect 1681 -1360 1685 -1340
rect 1725 -1360 1729 -1340
rect 1733 -1360 1737 -1340
rect 1773 -1343 1777 -1323
rect 1781 -1343 1785 -1323
rect 1805 -1343 1809 -1323
rect 1813 -1343 1817 -1323
rect 253 -1368 257 -1362
rect 261 -1368 265 -1362
rect 174 -1376 178 -1371
rect 198 -1376 202 -1371
rect -237 -1479 -233 -1459
rect -229 -1479 -225 -1459
rect -185 -1479 -181 -1459
rect -177 -1479 -173 -1459
rect 1334 -1465 1338 -1459
rect 1342 -1465 1346 -1459
rect 1256 -1473 1260 -1468
rect 1280 -1473 1284 -1468
rect -341 -1526 -337 -1506
rect -333 -1526 -329 -1506
rect -289 -1526 -285 -1506
rect -281 -1526 -277 -1506
rect -237 -1526 -233 -1506
rect -229 -1526 -225 -1506
rect -185 -1526 -181 -1506
rect -177 -1526 -173 -1506
rect -137 -1509 -133 -1489
rect -129 -1509 -125 -1489
rect -105 -1509 -101 -1489
rect -97 -1509 -93 -1489
rect 1435 -1515 1439 -1509
rect 1443 -1515 1447 -1509
rect 1394 -1521 1398 -1515
rect 1403 -1521 1407 -1515
rect 1412 -1521 1416 -1515
rect 1334 -1570 1338 -1564
rect 1342 -1570 1346 -1564
rect 1256 -1578 1260 -1573
rect 1280 -1578 1284 -1573
rect 1548 -1628 1552 -1622
rect 1556 -1628 1560 -1622
rect 1507 -1634 1511 -1628
rect 1516 -1634 1520 -1628
rect 1525 -1634 1529 -1628
rect -235 -1705 -231 -1685
rect -227 -1705 -223 -1685
rect -183 -1705 -179 -1685
rect -175 -1705 -171 -1685
rect 1334 -1673 1338 -1667
rect 1342 -1673 1346 -1667
rect 1256 -1681 1260 -1676
rect 1280 -1681 1284 -1676
rect -339 -1752 -335 -1732
rect -331 -1752 -327 -1732
rect -287 -1752 -283 -1732
rect -279 -1752 -275 -1732
rect -235 -1752 -231 -1732
rect -227 -1752 -223 -1732
rect -183 -1752 -179 -1732
rect -175 -1752 -171 -1732
rect -135 -1735 -131 -1715
rect -127 -1735 -123 -1715
rect -103 -1735 -99 -1715
rect -95 -1735 -91 -1715
rect 1432 -1717 1436 -1711
rect 1440 -1717 1444 -1711
rect 1391 -1723 1395 -1717
rect 1400 -1723 1404 -1717
rect 1409 -1723 1413 -1717
rect 1651 -1730 1655 -1724
rect 1659 -1730 1663 -1724
rect 1610 -1736 1614 -1730
rect 1619 -1736 1623 -1730
rect 1628 -1736 1632 -1730
rect 1324 -1762 1328 -1756
rect 1332 -1762 1336 -1756
rect 1246 -1770 1250 -1765
rect 1270 -1770 1274 -1765
rect -235 -1928 -231 -1908
rect -227 -1928 -223 -1908
rect -183 -1928 -179 -1908
rect -175 -1928 -171 -1908
rect -339 -1975 -335 -1955
rect -331 -1975 -327 -1955
rect -287 -1975 -283 -1955
rect -279 -1975 -275 -1955
rect -235 -1975 -231 -1955
rect -227 -1975 -223 -1955
rect -183 -1975 -179 -1955
rect -175 -1975 -171 -1955
rect -135 -1958 -131 -1938
rect -127 -1958 -123 -1938
rect -103 -1958 -99 -1938
rect -95 -1958 -91 -1938
<< pdcontact >>
rect -326 -306 -322 -266
rect -318 -306 -314 -266
rect -274 -306 -270 -266
rect -266 -306 -262 -266
rect -222 -306 -218 -266
rect -214 -306 -210 -266
rect -170 -306 -166 -266
rect -162 -306 -158 -266
rect -326 -368 -322 -328
rect -318 -368 -314 -328
rect -274 -368 -270 -328
rect -266 -368 -262 -328
rect -122 -352 -118 -312
rect -114 -352 -110 -312
rect -90 -352 -86 -312
rect -82 -352 -78 -312
rect 1581 -320 1585 -280
rect 1589 -320 1593 -280
rect 1633 -320 1637 -280
rect 1641 -320 1645 -280
rect 1685 -320 1689 -280
rect 1693 -320 1697 -280
rect 1737 -320 1741 -280
rect 1745 -320 1749 -280
rect 1581 -382 1585 -342
rect 1589 -382 1593 -342
rect 1633 -382 1637 -342
rect 1641 -382 1645 -342
rect 1785 -366 1789 -326
rect 1793 -366 1797 -326
rect 1817 -366 1821 -326
rect 1825 -366 1829 -326
rect 150 -469 154 -461
rect 158 -469 162 -461
rect 180 -469 184 -461
rect 200 -469 204 -461
rect 220 -469 224 -461
rect -329 -533 -325 -493
rect -321 -533 -317 -493
rect -277 -533 -273 -493
rect -269 -533 -265 -493
rect -225 -533 -221 -493
rect -217 -533 -213 -493
rect -173 -533 -169 -493
rect -165 -533 -161 -493
rect 150 -519 154 -511
rect 158 -519 162 -511
rect -329 -595 -325 -555
rect -321 -595 -317 -555
rect -277 -595 -273 -555
rect -269 -595 -265 -555
rect -125 -579 -121 -539
rect -117 -579 -113 -539
rect -93 -579 -89 -539
rect -85 -579 -81 -539
rect 963 -539 967 -531
rect 971 -539 975 -531
rect 993 -539 997 -531
rect 1013 -539 1017 -531
rect 1033 -539 1037 -531
rect 151 -590 155 -582
rect 159 -590 163 -582
rect 181 -590 185 -582
rect 201 -590 205 -582
rect 221 -590 225 -582
rect 151 -640 155 -632
rect 159 -640 163 -632
rect 963 -589 967 -581
rect 971 -589 975 -581
rect 1573 -562 1577 -522
rect 1581 -562 1585 -522
rect 1625 -562 1629 -522
rect 1633 -562 1637 -522
rect 1677 -562 1681 -522
rect 1685 -562 1689 -522
rect 1729 -562 1733 -522
rect 1737 -562 1741 -522
rect 633 -633 637 -628
rect 645 -633 649 -628
rect 657 -633 661 -628
rect 715 -653 719 -641
rect 723 -653 727 -641
rect 784 -653 788 -629
rect 802 -653 806 -629
rect 1573 -624 1577 -584
rect 1581 -624 1585 -584
rect 1625 -624 1629 -584
rect 1633 -624 1637 -584
rect 1777 -608 1781 -568
rect 1785 -608 1789 -568
rect 1809 -608 1813 -568
rect 1817 -608 1821 -568
rect 825 -654 829 -642
rect 833 -654 837 -642
rect 973 -663 977 -655
rect 981 -663 985 -655
rect 1003 -663 1007 -655
rect 1023 -663 1027 -655
rect 1043 -663 1047 -655
rect 151 -711 155 -703
rect 159 -711 163 -703
rect 181 -711 185 -703
rect 201 -711 205 -703
rect 221 -711 225 -703
rect -332 -762 -328 -722
rect -324 -762 -320 -722
rect -280 -762 -276 -722
rect -272 -762 -268 -722
rect -228 -762 -224 -722
rect -220 -762 -216 -722
rect -176 -762 -172 -722
rect -168 -762 -164 -722
rect 151 -761 155 -753
rect 159 -761 163 -753
rect -332 -824 -328 -784
rect -324 -824 -320 -784
rect -280 -824 -276 -784
rect -272 -824 -268 -784
rect -128 -808 -124 -768
rect -120 -808 -116 -768
rect -96 -808 -92 -768
rect -88 -808 -84 -768
rect 973 -713 977 -705
rect 981 -713 985 -705
rect 496 -718 500 -714
rect 507 -739 511 -735
rect 516 -718 520 -714
rect 527 -739 531 -734
rect 554 -724 559 -717
rect 564 -737 569 -732
rect 607 -773 611 -749
rect 625 -773 629 -749
rect 648 -774 652 -762
rect 656 -774 660 -762
rect 1574 -798 1578 -758
rect 1582 -798 1586 -758
rect 1626 -798 1630 -758
rect 1634 -798 1638 -758
rect 1678 -798 1682 -758
rect 1686 -798 1690 -758
rect 1730 -798 1734 -758
rect 1738 -798 1742 -758
rect 151 -831 155 -823
rect 159 -831 163 -823
rect 181 -831 185 -823
rect 201 -831 205 -823
rect 221 -831 225 -823
rect 151 -881 155 -873
rect 159 -881 163 -873
rect 877 -817 881 -809
rect 885 -817 889 -809
rect 907 -817 911 -809
rect 927 -817 931 -809
rect 947 -817 951 -809
rect 494 -824 498 -819
rect 506 -824 510 -819
rect 518 -824 522 -819
rect 571 -844 575 -832
rect 579 -844 583 -832
rect 646 -881 650 -857
rect 664 -881 668 -857
rect 877 -867 881 -859
rect 885 -867 889 -859
rect 687 -882 691 -870
rect 695 -882 699 -870
rect 1574 -860 1578 -820
rect 1582 -860 1586 -820
rect 1626 -860 1630 -820
rect 1634 -860 1638 -820
rect 1778 -844 1782 -804
rect 1786 -844 1790 -804
rect 1810 -844 1814 -804
rect 1818 -844 1822 -804
rect -332 -978 -328 -938
rect -324 -978 -320 -938
rect -280 -978 -276 -938
rect -272 -978 -268 -938
rect -228 -978 -224 -938
rect -220 -978 -216 -938
rect -176 -978 -172 -938
rect -168 -978 -164 -938
rect -332 -1040 -328 -1000
rect -324 -1040 -320 -1000
rect -280 -1040 -276 -1000
rect -272 -1040 -268 -1000
rect -128 -1024 -124 -984
rect -120 -1024 -116 -984
rect -96 -1024 -92 -984
rect -88 -1024 -84 -984
rect 852 -994 856 -989
rect 864 -994 868 -989
rect 876 -994 880 -989
rect 930 -1014 934 -1002
rect 938 -1014 942 -1002
rect 1574 -1031 1578 -991
rect 1582 -1031 1586 -991
rect 1626 -1031 1630 -991
rect 1634 -1031 1638 -991
rect 1678 -1031 1682 -991
rect 1686 -1031 1690 -991
rect 1730 -1031 1734 -991
rect 1738 -1031 1742 -991
rect 171 -1067 175 -1062
rect 183 -1067 187 -1062
rect 195 -1067 199 -1062
rect 249 -1087 253 -1075
rect 257 -1087 261 -1075
rect 1006 -1076 1010 -1052
rect 1024 -1076 1028 -1052
rect 856 -1101 860 -1096
rect 868 -1101 872 -1096
rect 880 -1101 884 -1096
rect 1047 -1077 1051 -1065
rect 1055 -1077 1059 -1065
rect 1321 -1103 1325 -1095
rect 1329 -1103 1333 -1095
rect 1351 -1103 1355 -1095
rect 1371 -1103 1375 -1095
rect 1391 -1103 1395 -1095
rect 934 -1121 938 -1109
rect 942 -1121 946 -1109
rect -333 -1193 -329 -1153
rect -325 -1193 -321 -1153
rect -281 -1193 -277 -1153
rect -273 -1193 -269 -1153
rect -229 -1193 -225 -1153
rect -221 -1193 -217 -1153
rect -177 -1193 -173 -1153
rect -169 -1193 -165 -1153
rect 172 -1154 176 -1149
rect 184 -1154 188 -1149
rect 196 -1154 200 -1149
rect 1094 -1155 1098 -1131
rect 1112 -1155 1116 -1131
rect 249 -1174 253 -1162
rect 257 -1174 261 -1162
rect 1135 -1156 1139 -1144
rect 1143 -1156 1147 -1144
rect 1321 -1153 1325 -1145
rect 1329 -1153 1333 -1145
rect 1574 -1093 1578 -1053
rect 1582 -1093 1586 -1053
rect 1626 -1093 1630 -1053
rect 1634 -1093 1638 -1053
rect 1778 -1077 1782 -1037
rect 1786 -1077 1790 -1037
rect 1810 -1077 1814 -1037
rect 1818 -1077 1822 -1037
rect -333 -1255 -329 -1215
rect -325 -1255 -321 -1215
rect -281 -1255 -277 -1215
rect -273 -1255 -269 -1215
rect -129 -1239 -125 -1199
rect -121 -1239 -117 -1199
rect -97 -1239 -93 -1199
rect -89 -1239 -85 -1199
rect 856 -1210 860 -1205
rect 868 -1210 872 -1205
rect 880 -1210 884 -1205
rect 174 -1242 178 -1237
rect 186 -1242 190 -1237
rect 198 -1242 202 -1237
rect 252 -1262 256 -1250
rect 260 -1262 264 -1250
rect 934 -1230 938 -1218
rect 942 -1230 946 -1218
rect 1006 -1245 1010 -1221
rect 1024 -1245 1028 -1221
rect 1047 -1246 1051 -1234
rect 1055 -1246 1059 -1234
rect 1569 -1257 1573 -1217
rect 1577 -1257 1581 -1217
rect 1621 -1257 1625 -1217
rect 1629 -1257 1633 -1217
rect 1673 -1257 1677 -1217
rect 1681 -1257 1685 -1217
rect 1725 -1257 1729 -1217
rect 1733 -1257 1737 -1217
rect 1569 -1319 1573 -1279
rect 1577 -1319 1581 -1279
rect 1621 -1319 1625 -1279
rect 1629 -1319 1633 -1279
rect 1773 -1303 1777 -1263
rect 1781 -1303 1785 -1263
rect 1805 -1303 1809 -1263
rect 1813 -1303 1817 -1263
rect 174 -1328 178 -1323
rect 186 -1328 190 -1323
rect 198 -1328 202 -1323
rect 253 -1348 257 -1336
rect 261 -1348 265 -1336
rect -341 -1423 -337 -1383
rect -333 -1423 -329 -1383
rect -289 -1423 -285 -1383
rect -281 -1423 -277 -1383
rect -237 -1423 -233 -1383
rect -229 -1423 -225 -1383
rect -185 -1423 -181 -1383
rect -177 -1423 -173 -1383
rect 1256 -1425 1260 -1420
rect -341 -1485 -337 -1445
rect -333 -1485 -329 -1445
rect -289 -1485 -285 -1445
rect -281 -1485 -277 -1445
rect -137 -1469 -133 -1429
rect -129 -1469 -125 -1429
rect -105 -1469 -101 -1429
rect -97 -1469 -93 -1429
rect 1268 -1425 1272 -1420
rect 1280 -1425 1284 -1420
rect 1334 -1445 1338 -1433
rect 1342 -1445 1346 -1433
rect 1394 -1494 1398 -1470
rect 1412 -1494 1416 -1470
rect 1435 -1495 1439 -1483
rect 1443 -1495 1447 -1483
rect 1256 -1530 1260 -1525
rect 1268 -1530 1272 -1525
rect 1280 -1530 1284 -1525
rect 1334 -1550 1338 -1538
rect 1342 -1550 1346 -1538
rect 1507 -1607 1511 -1583
rect 1525 -1607 1529 -1583
rect -339 -1649 -335 -1609
rect -331 -1649 -327 -1609
rect -287 -1649 -283 -1609
rect -279 -1649 -275 -1609
rect -235 -1649 -231 -1609
rect -227 -1649 -223 -1609
rect -183 -1649 -179 -1609
rect -175 -1649 -171 -1609
rect 1548 -1608 1552 -1596
rect 1556 -1608 1560 -1596
rect 1256 -1633 1260 -1628
rect 1268 -1633 1272 -1628
rect 1280 -1633 1284 -1628
rect -339 -1711 -335 -1671
rect -331 -1711 -327 -1671
rect -287 -1711 -283 -1671
rect -279 -1711 -275 -1671
rect -135 -1695 -131 -1655
rect -127 -1695 -123 -1655
rect -103 -1695 -99 -1655
rect -95 -1695 -91 -1655
rect 1334 -1653 1338 -1641
rect 1342 -1653 1346 -1641
rect 1391 -1696 1395 -1672
rect 1409 -1696 1413 -1672
rect 1432 -1697 1436 -1685
rect 1440 -1697 1444 -1685
rect 1610 -1709 1614 -1685
rect 1628 -1709 1632 -1685
rect 1246 -1722 1250 -1717
rect 1258 -1722 1262 -1717
rect 1270 -1722 1274 -1717
rect 1651 -1710 1655 -1698
rect 1659 -1710 1663 -1698
rect 1324 -1742 1328 -1730
rect 1332 -1742 1336 -1730
rect -339 -1872 -335 -1832
rect -331 -1872 -327 -1832
rect -287 -1872 -283 -1832
rect -279 -1872 -275 -1832
rect -235 -1872 -231 -1832
rect -227 -1872 -223 -1832
rect -183 -1872 -179 -1832
rect -175 -1872 -171 -1832
rect -339 -1934 -335 -1894
rect -331 -1934 -327 -1894
rect -287 -1934 -283 -1894
rect -279 -1934 -275 -1894
rect -135 -1918 -131 -1878
rect -127 -1918 -123 -1878
rect -103 -1918 -99 -1878
rect -95 -1918 -91 -1878
<< psubstratepcontact >>
rect -130 -405 -126 -401
rect -106 -405 -102 -401
rect -98 -405 -94 -401
rect -74 -405 -70 -401
rect -309 -422 -305 -418
rect -257 -422 -253 -418
rect -205 -422 -201 -418
rect -153 -422 -149 -418
rect 1777 -419 1781 -415
rect 1801 -419 1805 -415
rect 1809 -419 1813 -415
rect 1833 -419 1837 -415
rect 1598 -436 1602 -432
rect 1650 -436 1654 -432
rect 1702 -436 1706 -432
rect 1754 -436 1758 -432
rect -133 -632 -129 -628
rect -109 -632 -105 -628
rect -101 -632 -97 -628
rect -77 -632 -73 -628
rect -312 -649 -308 -645
rect -260 -649 -256 -645
rect -208 -649 -204 -645
rect -156 -649 -152 -645
rect 1769 -661 1773 -657
rect 1793 -661 1797 -657
rect 1801 -661 1805 -657
rect 1825 -661 1829 -657
rect 1590 -678 1594 -674
rect 1642 -678 1646 -674
rect 1694 -678 1698 -674
rect 1746 -678 1750 -674
rect 549 -782 572 -777
rect 497 -794 501 -790
rect 505 -794 509 -790
rect 513 -794 517 -790
rect 521 -794 525 -790
rect -136 -861 -132 -857
rect -112 -861 -108 -857
rect -104 -861 -100 -857
rect -80 -861 -76 -857
rect -315 -878 -311 -874
rect -263 -878 -259 -874
rect -211 -878 -207 -874
rect -159 -878 -155 -874
rect 1770 -897 1774 -893
rect 1794 -897 1798 -893
rect 1802 -897 1806 -893
rect 1826 -897 1830 -893
rect 1591 -914 1595 -910
rect 1643 -914 1647 -910
rect 1695 -914 1699 -910
rect 1747 -914 1751 -910
rect -136 -1077 -132 -1073
rect -112 -1077 -108 -1073
rect -104 -1077 -100 -1073
rect -80 -1077 -76 -1073
rect -315 -1094 -311 -1090
rect -263 -1094 -259 -1090
rect -211 -1094 -207 -1090
rect -159 -1094 -155 -1090
rect 1770 -1130 1774 -1126
rect 1794 -1130 1798 -1126
rect 1802 -1130 1806 -1126
rect 1826 -1130 1830 -1126
rect 1591 -1147 1595 -1143
rect 1643 -1147 1647 -1143
rect 1695 -1147 1699 -1143
rect 1747 -1147 1751 -1143
rect -137 -1292 -133 -1288
rect -113 -1292 -109 -1288
rect -105 -1292 -101 -1288
rect -81 -1292 -77 -1288
rect -316 -1309 -312 -1305
rect -264 -1309 -260 -1305
rect -212 -1309 -208 -1305
rect -160 -1309 -156 -1305
rect 1765 -1356 1769 -1352
rect 1789 -1356 1793 -1352
rect 1797 -1356 1801 -1352
rect 1821 -1356 1825 -1352
rect 1586 -1373 1590 -1369
rect 1638 -1373 1642 -1369
rect 1690 -1373 1694 -1369
rect 1742 -1373 1746 -1369
rect -145 -1522 -141 -1518
rect -121 -1522 -117 -1518
rect -113 -1522 -109 -1518
rect -89 -1522 -85 -1518
rect -324 -1539 -320 -1535
rect -272 -1539 -268 -1535
rect -220 -1539 -216 -1535
rect -168 -1539 -164 -1535
rect -143 -1748 -139 -1744
rect -119 -1748 -115 -1744
rect -111 -1748 -107 -1744
rect -87 -1748 -83 -1744
rect -322 -1765 -318 -1761
rect -270 -1765 -266 -1761
rect -218 -1765 -214 -1761
rect -166 -1765 -162 -1761
rect -143 -1971 -139 -1967
rect -119 -1971 -115 -1967
rect -111 -1971 -107 -1967
rect -87 -1971 -83 -1967
rect -322 -1988 -318 -1984
rect -270 -1988 -266 -1984
rect -218 -1988 -214 -1984
rect -166 -1988 -162 -1984
<< nsubstratencontact >>
rect -333 -258 -329 -254
rect -311 -258 -307 -254
rect -281 -258 -277 -254
rect -259 -258 -255 -254
rect -229 -258 -225 -254
rect -207 -258 -203 -254
rect -177 -258 -173 -254
rect -155 -258 -151 -254
rect 1574 -272 1578 -268
rect 1596 -272 1600 -268
rect 1626 -272 1630 -268
rect 1648 -272 1652 -268
rect 1678 -272 1682 -268
rect 1700 -272 1704 -268
rect 1730 -272 1734 -268
rect 1752 -272 1756 -268
rect -129 -304 -125 -300
rect -107 -304 -103 -300
rect -97 -304 -93 -300
rect -75 -304 -71 -300
rect 1778 -318 1782 -314
rect 1800 -318 1804 -314
rect 1810 -318 1814 -314
rect 1832 -318 1836 -314
rect -336 -485 -332 -481
rect -314 -485 -310 -481
rect -284 -485 -280 -481
rect -262 -485 -258 -481
rect -232 -485 -228 -481
rect -210 -485 -206 -481
rect -180 -485 -176 -481
rect -158 -485 -154 -481
rect -132 -531 -128 -527
rect -110 -531 -106 -527
rect -100 -531 -96 -527
rect -78 -531 -74 -527
rect 1566 -514 1570 -510
rect 1588 -514 1592 -510
rect 1618 -514 1622 -510
rect 1640 -514 1644 -510
rect 1670 -514 1674 -510
rect 1692 -514 1696 -510
rect 1722 -514 1726 -510
rect 1744 -514 1748 -510
rect 1770 -560 1774 -556
rect 1792 -560 1796 -556
rect 1802 -560 1806 -556
rect 1824 -560 1828 -556
rect -339 -714 -335 -710
rect -317 -714 -313 -710
rect -287 -714 -283 -710
rect -265 -714 -261 -710
rect -235 -714 -231 -710
rect -213 -714 -209 -710
rect -183 -714 -179 -710
rect -161 -714 -157 -710
rect -135 -760 -131 -756
rect -113 -760 -109 -756
rect -103 -760 -99 -756
rect -81 -760 -77 -756
rect 497 -704 501 -700
rect 509 -704 513 -700
rect 518 -704 522 -700
rect 526 -704 530 -700
rect 550 -710 554 -706
rect 558 -710 562 -706
rect 566 -710 570 -706
rect 1567 -750 1571 -746
rect 1589 -750 1593 -746
rect 1619 -750 1623 -746
rect 1641 -750 1645 -746
rect 1671 -750 1675 -746
rect 1693 -750 1697 -746
rect 1723 -750 1727 -746
rect 1745 -750 1749 -746
rect 1771 -796 1775 -792
rect 1793 -796 1797 -792
rect 1803 -796 1807 -792
rect 1825 -796 1829 -792
rect -339 -930 -335 -926
rect -317 -930 -313 -926
rect -287 -930 -283 -926
rect -265 -930 -261 -926
rect -235 -930 -231 -926
rect -213 -930 -209 -926
rect -183 -930 -179 -926
rect -161 -930 -157 -926
rect -135 -976 -131 -972
rect -113 -976 -109 -972
rect -103 -976 -99 -972
rect -81 -976 -77 -972
rect 1567 -983 1571 -979
rect 1589 -983 1593 -979
rect 1619 -983 1623 -979
rect 1641 -983 1645 -979
rect 1671 -983 1675 -979
rect 1693 -983 1697 -979
rect 1723 -983 1727 -979
rect 1745 -983 1749 -979
rect 1771 -1029 1775 -1025
rect 1793 -1029 1797 -1025
rect 1803 -1029 1807 -1025
rect 1825 -1029 1829 -1025
rect -340 -1145 -336 -1141
rect -318 -1145 -314 -1141
rect -288 -1145 -284 -1141
rect -266 -1145 -262 -1141
rect -236 -1145 -232 -1141
rect -214 -1145 -210 -1141
rect -184 -1145 -180 -1141
rect -162 -1145 -158 -1141
rect -136 -1191 -132 -1187
rect -114 -1191 -110 -1187
rect -104 -1191 -100 -1187
rect -82 -1191 -78 -1187
rect 1562 -1209 1566 -1205
rect 1584 -1209 1588 -1205
rect 1614 -1209 1618 -1205
rect 1636 -1209 1640 -1205
rect 1666 -1209 1670 -1205
rect 1688 -1209 1692 -1205
rect 1718 -1209 1722 -1205
rect 1740 -1209 1744 -1205
rect 1766 -1255 1770 -1251
rect 1788 -1255 1792 -1251
rect 1798 -1255 1802 -1251
rect 1820 -1255 1824 -1251
rect -348 -1375 -344 -1371
rect -326 -1375 -322 -1371
rect -296 -1375 -292 -1371
rect -274 -1375 -270 -1371
rect -244 -1375 -240 -1371
rect -222 -1375 -218 -1371
rect -192 -1375 -188 -1371
rect -170 -1375 -166 -1371
rect -144 -1421 -140 -1417
rect -122 -1421 -118 -1417
rect -112 -1421 -108 -1417
rect -90 -1421 -86 -1417
rect -346 -1601 -342 -1597
rect -324 -1601 -320 -1597
rect -294 -1601 -290 -1597
rect -272 -1601 -268 -1597
rect -242 -1601 -238 -1597
rect -220 -1601 -216 -1597
rect -190 -1601 -186 -1597
rect -168 -1601 -164 -1597
rect -142 -1647 -138 -1643
rect -120 -1647 -116 -1643
rect -110 -1647 -106 -1643
rect -88 -1647 -84 -1643
rect -346 -1824 -342 -1820
rect -324 -1824 -320 -1820
rect -294 -1824 -290 -1820
rect -272 -1824 -268 -1820
rect -242 -1824 -238 -1820
rect -220 -1824 -216 -1820
rect -190 -1824 -186 -1820
rect -168 -1824 -164 -1820
rect -142 -1870 -138 -1866
rect -120 -1870 -116 -1866
rect -110 -1870 -106 -1866
rect -88 -1870 -84 -1866
<< polysilicon >>
rect -321 -266 -319 -262
rect -269 -266 -267 -262
rect -217 -266 -215 -262
rect -165 -266 -163 -262
rect 1586 -280 1588 -276
rect 1638 -280 1640 -276
rect 1690 -280 1692 -276
rect 1742 -280 1744 -276
rect -321 -315 -319 -306
rect -269 -315 -267 -306
rect -217 -315 -215 -306
rect -165 -315 -163 -306
rect -117 -312 -115 -308
rect -85 -312 -83 -308
rect -321 -328 -319 -324
rect -269 -328 -267 -324
rect -217 -342 -215 -333
rect -165 -342 -163 -333
rect 1586 -329 1588 -320
rect 1638 -329 1640 -320
rect 1690 -329 1692 -320
rect 1742 -329 1744 -320
rect 1790 -326 1792 -322
rect 1822 -326 1824 -322
rect 1586 -342 1588 -338
rect 1638 -342 1640 -338
rect -217 -365 -215 -362
rect -165 -365 -163 -362
rect -321 -377 -319 -368
rect -269 -377 -267 -368
rect -117 -372 -115 -352
rect -85 -372 -83 -352
rect -321 -389 -319 -381
rect -269 -389 -267 -381
rect -217 -389 -215 -381
rect -165 -389 -163 -381
rect 1690 -356 1692 -347
rect 1742 -356 1744 -347
rect 1690 -379 1692 -376
rect 1742 -379 1744 -376
rect 1586 -391 1588 -382
rect 1638 -391 1640 -382
rect 1790 -386 1792 -366
rect 1822 -386 1824 -366
rect -117 -396 -115 -392
rect -85 -396 -83 -392
rect 1586 -403 1588 -395
rect 1638 -403 1640 -395
rect 1690 -403 1692 -395
rect 1742 -403 1744 -395
rect -321 -413 -319 -409
rect -269 -413 -267 -409
rect -217 -413 -215 -409
rect -165 -413 -163 -409
rect 1790 -410 1792 -406
rect 1822 -410 1824 -406
rect 1586 -427 1588 -423
rect 1638 -427 1640 -423
rect 1690 -427 1692 -423
rect 1742 -427 1744 -423
rect 186 -451 228 -449
rect 155 -461 157 -458
rect 186 -461 188 -451
rect 196 -461 198 -458
rect 206 -461 208 -458
rect 216 -461 218 -458
rect 155 -483 157 -469
rect 186 -480 188 -469
rect 196 -484 198 -469
rect 186 -486 198 -484
rect -324 -493 -322 -489
rect -272 -493 -270 -489
rect -220 -493 -218 -489
rect -168 -493 -166 -489
rect 155 -490 157 -487
rect 155 -511 157 -508
rect 155 -533 157 -519
rect 186 -533 188 -486
rect 206 -489 208 -469
rect 196 -491 208 -489
rect 196 -533 198 -491
rect 216 -523 218 -469
rect 206 -525 218 -523
rect 206 -533 208 -525
rect 226 -528 228 -451
rect 999 -521 1041 -519
rect 216 -530 228 -528
rect 216 -533 218 -530
rect 968 -531 970 -528
rect 999 -531 1001 -521
rect 1009 -531 1011 -528
rect 1019 -531 1021 -528
rect 1029 -531 1031 -528
rect -324 -542 -322 -533
rect -272 -542 -270 -533
rect -220 -542 -218 -533
rect -168 -542 -166 -533
rect -120 -539 -118 -535
rect -88 -539 -86 -535
rect -324 -555 -322 -551
rect -272 -555 -270 -551
rect -220 -569 -218 -560
rect -168 -569 -166 -560
rect 155 -540 157 -537
rect 186 -553 188 -537
rect 196 -540 198 -537
rect 206 -561 208 -537
rect 216 -540 218 -537
rect 968 -553 970 -539
rect 999 -550 1001 -539
rect 1009 -554 1011 -539
rect 999 -556 1011 -554
rect 968 -560 970 -557
rect 187 -572 229 -570
rect -220 -592 -218 -589
rect -168 -592 -166 -589
rect -324 -604 -322 -595
rect -272 -604 -270 -595
rect -120 -599 -118 -579
rect -88 -599 -86 -579
rect 156 -582 158 -579
rect 187 -582 189 -572
rect 197 -582 199 -579
rect 207 -582 209 -579
rect 217 -582 219 -579
rect -324 -616 -322 -608
rect -272 -616 -270 -608
rect -220 -616 -218 -608
rect -168 -616 -166 -608
rect 156 -604 158 -590
rect 187 -601 189 -590
rect 197 -605 199 -590
rect 187 -607 199 -605
rect 156 -611 158 -608
rect -120 -623 -118 -619
rect -88 -623 -86 -619
rect 156 -632 158 -629
rect -324 -640 -322 -636
rect -272 -640 -270 -636
rect -220 -640 -218 -636
rect -168 -640 -166 -636
rect 156 -654 158 -640
rect 187 -654 189 -607
rect 207 -610 209 -590
rect 197 -612 209 -610
rect 197 -654 199 -612
rect 217 -644 219 -590
rect 207 -646 219 -644
rect 207 -654 209 -646
rect 227 -649 229 -572
rect 968 -581 970 -578
rect 968 -603 970 -589
rect 999 -603 1001 -556
rect 1019 -559 1021 -539
rect 1009 -561 1021 -559
rect 1009 -603 1011 -561
rect 1029 -593 1031 -539
rect 1019 -595 1031 -593
rect 1019 -603 1021 -595
rect 1039 -598 1041 -521
rect 1578 -522 1580 -518
rect 1630 -522 1632 -518
rect 1682 -522 1684 -518
rect 1734 -522 1736 -518
rect 1578 -571 1580 -562
rect 1630 -571 1632 -562
rect 1682 -571 1684 -562
rect 1734 -571 1736 -562
rect 1782 -568 1784 -564
rect 1814 -568 1816 -564
rect 1578 -584 1580 -580
rect 1630 -584 1632 -580
rect 1029 -600 1041 -598
rect 1029 -603 1031 -600
rect 968 -610 970 -607
rect 999 -623 1001 -607
rect 1009 -610 1011 -607
rect 639 -628 642 -624
rect 652 -628 655 -624
rect 789 -629 791 -626
rect 799 -629 801 -626
rect 720 -641 722 -638
rect 217 -651 229 -649
rect 217 -654 219 -651
rect 639 -657 642 -648
rect 156 -661 158 -658
rect 187 -674 189 -658
rect 197 -661 199 -658
rect 207 -682 209 -658
rect 217 -661 219 -658
rect 641 -661 642 -657
rect 639 -676 642 -661
rect 652 -668 655 -648
rect 1019 -631 1021 -607
rect 1029 -610 1031 -607
rect 1682 -598 1684 -589
rect 1734 -598 1736 -589
rect 1682 -621 1684 -618
rect 1734 -621 1736 -618
rect 1578 -633 1580 -624
rect 1630 -633 1632 -624
rect 1782 -628 1784 -608
rect 1814 -628 1816 -608
rect 830 -642 832 -639
rect 720 -667 722 -653
rect 654 -672 655 -668
rect 652 -676 655 -672
rect 720 -676 722 -673
rect 789 -674 791 -653
rect 799 -674 801 -653
rect 1009 -645 1051 -643
rect 1578 -645 1580 -637
rect 1630 -645 1632 -637
rect 1682 -645 1684 -637
rect 1734 -645 1736 -637
rect 830 -668 832 -654
rect 978 -655 980 -652
rect 1009 -655 1011 -645
rect 1019 -655 1021 -652
rect 1029 -655 1031 -652
rect 1039 -655 1041 -652
rect 187 -693 229 -691
rect 830 -677 832 -674
rect 978 -677 980 -663
rect 1009 -674 1011 -663
rect 789 -683 791 -680
rect 799 -683 801 -680
rect 1019 -678 1021 -663
rect 1009 -680 1021 -678
rect 978 -684 980 -681
rect 156 -703 158 -700
rect 187 -703 189 -693
rect 197 -703 199 -700
rect 207 -703 209 -700
rect 217 -703 219 -700
rect -327 -722 -325 -718
rect -275 -722 -273 -718
rect -223 -722 -221 -718
rect -171 -722 -169 -718
rect 156 -725 158 -711
rect 187 -722 189 -711
rect 197 -726 199 -711
rect 187 -728 199 -726
rect 156 -732 158 -729
rect 156 -753 158 -750
rect -327 -771 -325 -762
rect -275 -771 -273 -762
rect -223 -771 -221 -762
rect -171 -771 -169 -762
rect -123 -768 -121 -764
rect -91 -768 -89 -764
rect -327 -784 -325 -780
rect -275 -784 -273 -780
rect -223 -798 -221 -789
rect -171 -798 -169 -789
rect 156 -775 158 -761
rect 187 -775 189 -728
rect 207 -731 209 -711
rect 197 -733 209 -731
rect 197 -775 199 -733
rect 217 -765 219 -711
rect 207 -767 219 -765
rect 207 -775 209 -767
rect 227 -770 229 -693
rect 639 -697 642 -692
rect 652 -697 655 -692
rect 978 -705 980 -702
rect 503 -714 505 -711
rect 513 -714 515 -711
rect 521 -714 523 -711
rect 560 -717 562 -713
rect 978 -727 980 -713
rect 1009 -727 1011 -680
rect 1029 -683 1031 -663
rect 1019 -685 1031 -683
rect 1019 -727 1021 -685
rect 1039 -717 1041 -663
rect 1029 -719 1041 -717
rect 1029 -727 1031 -719
rect 1049 -722 1051 -645
rect 1782 -652 1784 -648
rect 1814 -652 1816 -648
rect 1578 -669 1580 -665
rect 1630 -669 1632 -665
rect 1682 -669 1684 -665
rect 1734 -669 1736 -665
rect 1039 -724 1051 -722
rect 1039 -727 1041 -724
rect 978 -734 980 -731
rect 503 -748 505 -739
rect 504 -754 505 -748
rect 217 -772 229 -770
rect 503 -771 505 -754
rect 513 -757 515 -739
rect 513 -771 515 -761
rect 521 -764 523 -739
rect 560 -749 562 -737
rect 612 -749 614 -746
rect 622 -749 624 -746
rect 1009 -747 1011 -731
rect 1019 -734 1021 -731
rect 561 -754 562 -749
rect 560 -758 562 -754
rect 521 -771 523 -768
rect 217 -775 219 -772
rect 156 -782 158 -779
rect 187 -795 189 -779
rect 197 -782 199 -779
rect 207 -803 209 -779
rect 217 -782 219 -779
rect 560 -773 562 -768
rect 1029 -755 1031 -731
rect 1039 -734 1041 -731
rect 1579 -758 1581 -754
rect 1631 -758 1633 -754
rect 1683 -758 1685 -754
rect 1735 -758 1737 -754
rect 653 -762 655 -759
rect 503 -785 505 -781
rect 513 -785 515 -781
rect 521 -786 523 -781
rect 612 -794 614 -773
rect 622 -794 624 -773
rect 653 -788 655 -774
rect 653 -797 655 -794
rect 913 -799 955 -797
rect 612 -803 614 -800
rect 622 -803 624 -800
rect -223 -821 -221 -818
rect -171 -821 -169 -818
rect -327 -833 -325 -824
rect -275 -833 -273 -824
rect -123 -828 -121 -808
rect -91 -828 -89 -808
rect 882 -809 884 -806
rect 913 -809 915 -799
rect 923 -809 925 -806
rect 933 -809 935 -806
rect 943 -809 945 -806
rect 187 -813 229 -811
rect 156 -823 158 -820
rect 187 -823 189 -813
rect 197 -823 199 -820
rect 207 -823 209 -820
rect 217 -823 219 -820
rect -327 -845 -325 -837
rect -275 -845 -273 -837
rect -223 -845 -221 -837
rect -171 -845 -169 -837
rect 156 -845 158 -831
rect 187 -842 189 -831
rect -123 -852 -121 -848
rect -91 -852 -89 -848
rect 197 -846 199 -831
rect 187 -848 199 -846
rect 156 -852 158 -849
rect -327 -869 -325 -865
rect -275 -869 -273 -865
rect -223 -869 -221 -865
rect -171 -869 -169 -865
rect 156 -873 158 -870
rect 156 -895 158 -881
rect 187 -895 189 -848
rect 207 -851 209 -831
rect 197 -853 209 -851
rect 197 -895 199 -853
rect 217 -885 219 -831
rect 207 -887 219 -885
rect 207 -895 209 -887
rect 227 -890 229 -813
rect 500 -819 503 -815
rect 513 -819 516 -815
rect 576 -832 578 -829
rect 882 -831 884 -817
rect 913 -828 915 -817
rect 500 -848 503 -839
rect 502 -852 503 -848
rect 500 -867 503 -852
rect 513 -859 516 -839
rect 923 -832 925 -817
rect 913 -834 925 -832
rect 882 -838 884 -835
rect 576 -858 578 -844
rect 651 -857 653 -854
rect 661 -857 663 -854
rect 515 -863 516 -859
rect 513 -867 516 -863
rect 576 -867 578 -864
rect 882 -859 884 -856
rect 692 -870 694 -867
rect 500 -888 503 -883
rect 513 -888 516 -883
rect 217 -892 229 -890
rect 217 -895 219 -892
rect 156 -902 158 -899
rect 187 -915 189 -899
rect 197 -902 199 -899
rect 207 -923 209 -899
rect 217 -902 219 -899
rect 651 -902 653 -881
rect 661 -902 663 -881
rect 882 -881 884 -867
rect 913 -881 915 -834
rect 933 -837 935 -817
rect 923 -839 935 -837
rect 923 -881 925 -839
rect 943 -871 945 -817
rect 933 -873 945 -871
rect 933 -881 935 -873
rect 953 -876 955 -799
rect 1579 -807 1581 -798
rect 1631 -807 1633 -798
rect 1683 -807 1685 -798
rect 1735 -807 1737 -798
rect 1783 -804 1785 -800
rect 1815 -804 1817 -800
rect 1579 -820 1581 -816
rect 1631 -820 1633 -816
rect 1683 -834 1685 -825
rect 1735 -834 1737 -825
rect 1683 -857 1685 -854
rect 1735 -857 1737 -854
rect 1579 -869 1581 -860
rect 1631 -869 1633 -860
rect 1783 -864 1785 -844
rect 1815 -864 1817 -844
rect 943 -878 955 -876
rect 943 -881 945 -878
rect 1579 -881 1581 -873
rect 1631 -881 1633 -873
rect 1683 -881 1685 -873
rect 1735 -881 1737 -873
rect 692 -896 694 -882
rect 882 -888 884 -885
rect 913 -901 915 -885
rect 923 -888 925 -885
rect 692 -905 694 -902
rect 651 -911 653 -908
rect 661 -911 663 -908
rect 933 -909 935 -885
rect 943 -888 945 -885
rect 1783 -888 1785 -884
rect 1815 -888 1817 -884
rect 1579 -905 1581 -901
rect 1631 -905 1633 -901
rect 1683 -905 1685 -901
rect 1735 -905 1737 -901
rect -327 -938 -325 -934
rect -275 -938 -273 -934
rect -223 -938 -221 -934
rect -171 -938 -169 -934
rect -327 -987 -325 -978
rect -275 -987 -273 -978
rect -223 -987 -221 -978
rect -171 -987 -169 -978
rect -123 -984 -121 -980
rect -91 -984 -89 -980
rect -327 -1000 -325 -996
rect -275 -1000 -273 -996
rect -223 -1014 -221 -1005
rect -171 -1014 -169 -1005
rect 858 -989 861 -985
rect 871 -989 874 -985
rect 1579 -991 1581 -987
rect 1631 -991 1633 -987
rect 1683 -991 1685 -987
rect 1735 -991 1737 -987
rect 935 -1002 937 -999
rect 858 -1018 861 -1009
rect 860 -1022 861 -1018
rect -223 -1037 -221 -1034
rect -171 -1037 -169 -1034
rect -327 -1049 -325 -1040
rect -275 -1049 -273 -1040
rect -123 -1044 -121 -1024
rect -91 -1044 -89 -1024
rect 858 -1037 861 -1022
rect 871 -1029 874 -1009
rect 935 -1028 937 -1014
rect 873 -1033 874 -1029
rect 871 -1037 874 -1033
rect 935 -1037 937 -1034
rect -327 -1061 -325 -1053
rect -275 -1061 -273 -1053
rect -223 -1061 -221 -1053
rect -171 -1061 -169 -1053
rect 1579 -1040 1581 -1031
rect 1631 -1040 1633 -1031
rect 1683 -1040 1685 -1031
rect 1735 -1040 1737 -1031
rect 1783 -1037 1785 -1033
rect 1815 -1037 1817 -1033
rect 1011 -1052 1013 -1049
rect 1021 -1052 1023 -1049
rect 858 -1058 861 -1053
rect 871 -1058 874 -1053
rect 177 -1062 180 -1058
rect 190 -1062 193 -1058
rect -123 -1068 -121 -1064
rect -91 -1068 -89 -1064
rect -327 -1085 -325 -1081
rect -275 -1085 -273 -1081
rect -223 -1085 -221 -1081
rect -171 -1085 -169 -1081
rect 254 -1075 256 -1072
rect 177 -1091 180 -1082
rect 179 -1095 180 -1091
rect 177 -1110 180 -1095
rect 190 -1102 193 -1082
rect 1579 -1053 1581 -1049
rect 1631 -1053 1633 -1049
rect 1052 -1065 1054 -1062
rect 254 -1101 256 -1087
rect 862 -1096 865 -1092
rect 875 -1096 878 -1092
rect 192 -1106 193 -1102
rect 190 -1110 193 -1106
rect 254 -1110 256 -1107
rect 1011 -1097 1013 -1076
rect 1021 -1097 1023 -1076
rect 1052 -1091 1054 -1077
rect 1357 -1085 1399 -1083
rect 1326 -1095 1328 -1092
rect 1357 -1095 1359 -1085
rect 1367 -1095 1369 -1092
rect 1377 -1095 1379 -1092
rect 1387 -1095 1389 -1092
rect 1052 -1100 1054 -1097
rect 1011 -1106 1013 -1103
rect 1021 -1106 1023 -1103
rect 939 -1109 941 -1106
rect 862 -1125 865 -1116
rect 177 -1131 180 -1126
rect 190 -1131 193 -1126
rect 864 -1129 865 -1125
rect 862 -1144 865 -1129
rect 875 -1136 878 -1116
rect 1326 -1117 1328 -1103
rect 1357 -1114 1359 -1103
rect 1367 -1118 1369 -1103
rect 1357 -1120 1369 -1118
rect 939 -1135 941 -1121
rect 1326 -1124 1328 -1121
rect 1099 -1131 1101 -1128
rect 1109 -1131 1111 -1128
rect 877 -1140 878 -1136
rect 875 -1144 878 -1140
rect 939 -1144 941 -1141
rect 178 -1149 181 -1145
rect 191 -1149 194 -1145
rect -328 -1153 -326 -1149
rect -276 -1153 -274 -1149
rect -224 -1153 -222 -1149
rect -172 -1153 -170 -1149
rect 254 -1162 256 -1159
rect 1140 -1144 1142 -1141
rect 178 -1178 181 -1169
rect 180 -1182 181 -1178
rect -328 -1202 -326 -1193
rect -276 -1202 -274 -1193
rect -224 -1202 -222 -1193
rect -172 -1202 -170 -1193
rect -124 -1199 -122 -1195
rect -92 -1199 -90 -1195
rect 178 -1197 181 -1182
rect 191 -1189 194 -1169
rect 862 -1165 865 -1160
rect 875 -1165 878 -1160
rect 254 -1188 256 -1174
rect 1099 -1176 1101 -1155
rect 1109 -1176 1111 -1155
rect 1326 -1145 1328 -1142
rect 1140 -1170 1142 -1156
rect 1326 -1167 1328 -1153
rect 1357 -1167 1359 -1120
rect 1377 -1123 1379 -1103
rect 1367 -1125 1379 -1123
rect 1367 -1167 1369 -1125
rect 1387 -1157 1389 -1103
rect 1377 -1159 1389 -1157
rect 1377 -1167 1379 -1159
rect 1397 -1162 1399 -1085
rect 1683 -1067 1685 -1058
rect 1735 -1067 1737 -1058
rect 1683 -1090 1685 -1087
rect 1735 -1090 1737 -1087
rect 1579 -1102 1581 -1093
rect 1631 -1102 1633 -1093
rect 1783 -1097 1785 -1077
rect 1815 -1097 1817 -1077
rect 1579 -1114 1581 -1106
rect 1631 -1114 1633 -1106
rect 1683 -1114 1685 -1106
rect 1735 -1114 1737 -1106
rect 1783 -1121 1785 -1117
rect 1815 -1121 1817 -1117
rect 1579 -1138 1581 -1134
rect 1631 -1138 1633 -1134
rect 1683 -1138 1685 -1134
rect 1735 -1138 1737 -1134
rect 1387 -1164 1399 -1162
rect 1387 -1167 1389 -1164
rect 1326 -1174 1328 -1171
rect 1140 -1179 1142 -1176
rect 1099 -1185 1101 -1182
rect 1109 -1185 1111 -1182
rect 1357 -1187 1359 -1171
rect 1367 -1174 1369 -1171
rect 193 -1193 194 -1189
rect 191 -1197 194 -1193
rect 254 -1197 256 -1194
rect 1377 -1195 1379 -1171
rect 1387 -1174 1389 -1171
rect -328 -1215 -326 -1211
rect -276 -1215 -274 -1211
rect -224 -1229 -222 -1220
rect -172 -1229 -170 -1220
rect 862 -1205 865 -1201
rect 875 -1205 878 -1201
rect 178 -1218 181 -1213
rect 191 -1218 194 -1213
rect 939 -1218 941 -1215
rect 1574 -1217 1576 -1213
rect 1626 -1217 1628 -1213
rect 1678 -1217 1680 -1213
rect 1730 -1217 1732 -1213
rect 180 -1237 183 -1233
rect 193 -1237 196 -1233
rect 862 -1234 865 -1225
rect -224 -1252 -222 -1249
rect -172 -1252 -170 -1249
rect -328 -1264 -326 -1255
rect -276 -1264 -274 -1255
rect -124 -1259 -122 -1239
rect -92 -1259 -90 -1239
rect 864 -1238 865 -1234
rect 257 -1250 259 -1247
rect -328 -1276 -326 -1268
rect -276 -1276 -274 -1268
rect -224 -1276 -222 -1268
rect -172 -1276 -170 -1268
rect 180 -1266 183 -1257
rect 182 -1270 183 -1266
rect -124 -1283 -122 -1279
rect -92 -1283 -90 -1279
rect 180 -1285 183 -1270
rect 193 -1277 196 -1257
rect 862 -1253 865 -1238
rect 875 -1245 878 -1225
rect 1011 -1221 1013 -1218
rect 1021 -1221 1023 -1218
rect 939 -1244 941 -1230
rect 877 -1249 878 -1245
rect 875 -1253 878 -1249
rect 1052 -1234 1054 -1231
rect 939 -1253 941 -1250
rect 257 -1276 259 -1262
rect 1011 -1266 1013 -1245
rect 1021 -1266 1023 -1245
rect 1052 -1260 1054 -1246
rect 1574 -1266 1576 -1257
rect 1626 -1266 1628 -1257
rect 1678 -1266 1680 -1257
rect 1730 -1266 1732 -1257
rect 1778 -1263 1780 -1259
rect 1810 -1263 1812 -1259
rect 862 -1274 865 -1269
rect 875 -1274 878 -1269
rect 1052 -1269 1054 -1266
rect 1011 -1275 1013 -1272
rect 1021 -1275 1023 -1272
rect 195 -1281 196 -1277
rect 193 -1285 196 -1281
rect 1574 -1279 1576 -1275
rect 1626 -1279 1628 -1275
rect 257 -1285 259 -1282
rect -328 -1300 -326 -1296
rect -276 -1300 -274 -1296
rect -224 -1300 -222 -1296
rect -172 -1300 -170 -1296
rect 180 -1306 183 -1301
rect 193 -1306 196 -1301
rect 1678 -1293 1680 -1284
rect 1730 -1293 1732 -1284
rect 1678 -1316 1680 -1313
rect 1730 -1316 1732 -1313
rect 180 -1323 183 -1319
rect 193 -1323 196 -1319
rect 1574 -1328 1576 -1319
rect 1626 -1328 1628 -1319
rect 1778 -1323 1780 -1303
rect 1810 -1323 1812 -1303
rect 258 -1336 260 -1333
rect 180 -1352 183 -1343
rect 182 -1356 183 -1352
rect 180 -1371 183 -1356
rect 193 -1363 196 -1343
rect 1574 -1340 1576 -1332
rect 1626 -1340 1628 -1332
rect 1678 -1340 1680 -1332
rect 1730 -1340 1732 -1332
rect 258 -1362 260 -1348
rect 1778 -1347 1780 -1343
rect 1810 -1347 1812 -1343
rect 195 -1367 196 -1363
rect 193 -1371 196 -1367
rect 1574 -1364 1576 -1360
rect 1626 -1364 1628 -1360
rect 1678 -1364 1680 -1360
rect 1730 -1364 1732 -1360
rect 258 -1371 260 -1368
rect -336 -1383 -334 -1379
rect -284 -1383 -282 -1379
rect -232 -1383 -230 -1379
rect -180 -1383 -178 -1379
rect 180 -1392 183 -1387
rect 193 -1392 196 -1387
rect 1262 -1420 1265 -1416
rect 1275 -1420 1278 -1416
rect -336 -1432 -334 -1423
rect -284 -1432 -282 -1423
rect -232 -1432 -230 -1423
rect -180 -1432 -178 -1423
rect -132 -1429 -130 -1425
rect -100 -1429 -98 -1425
rect -336 -1445 -334 -1441
rect -284 -1445 -282 -1441
rect -232 -1459 -230 -1450
rect -180 -1459 -178 -1450
rect 1339 -1433 1341 -1430
rect 1262 -1449 1265 -1440
rect 1264 -1453 1265 -1449
rect 1262 -1468 1265 -1453
rect 1275 -1460 1278 -1440
rect 1339 -1459 1341 -1445
rect 1277 -1464 1278 -1460
rect 1275 -1468 1278 -1464
rect 1339 -1468 1341 -1465
rect -232 -1482 -230 -1479
rect -180 -1482 -178 -1479
rect -336 -1494 -334 -1485
rect -284 -1494 -282 -1485
rect -132 -1489 -130 -1469
rect -100 -1489 -98 -1469
rect 1399 -1470 1401 -1467
rect 1409 -1470 1411 -1467
rect 1262 -1489 1265 -1484
rect 1275 -1489 1278 -1484
rect -336 -1506 -334 -1498
rect -284 -1506 -282 -1498
rect -232 -1506 -230 -1498
rect -180 -1506 -178 -1498
rect 1440 -1483 1442 -1480
rect -132 -1513 -130 -1509
rect -100 -1513 -98 -1509
rect 1399 -1515 1401 -1494
rect 1409 -1515 1411 -1494
rect 1440 -1509 1442 -1495
rect 1440 -1518 1442 -1515
rect 1262 -1525 1265 -1521
rect 1275 -1525 1278 -1521
rect 1399 -1524 1401 -1521
rect 1409 -1524 1411 -1521
rect -336 -1530 -334 -1526
rect -284 -1530 -282 -1526
rect -232 -1530 -230 -1526
rect -180 -1530 -178 -1526
rect 1339 -1538 1341 -1535
rect 1262 -1554 1265 -1545
rect 1264 -1558 1265 -1554
rect 1262 -1573 1265 -1558
rect 1275 -1565 1278 -1545
rect 1339 -1564 1341 -1550
rect 1277 -1569 1278 -1565
rect 1275 -1573 1278 -1569
rect 1339 -1573 1341 -1570
rect 1512 -1583 1514 -1580
rect 1522 -1583 1524 -1580
rect 1262 -1594 1265 -1589
rect 1275 -1594 1278 -1589
rect -334 -1609 -332 -1605
rect -282 -1609 -280 -1605
rect -230 -1609 -228 -1605
rect -178 -1609 -176 -1605
rect 1553 -1596 1555 -1593
rect 1262 -1628 1265 -1624
rect 1275 -1628 1278 -1624
rect 1512 -1628 1514 -1607
rect 1522 -1628 1524 -1607
rect 1553 -1622 1555 -1608
rect 1553 -1631 1555 -1628
rect 1512 -1637 1514 -1634
rect 1522 -1637 1524 -1634
rect 1339 -1641 1341 -1638
rect -334 -1658 -332 -1649
rect -282 -1658 -280 -1649
rect -230 -1658 -228 -1649
rect -178 -1658 -176 -1649
rect -130 -1655 -128 -1651
rect -98 -1655 -96 -1651
rect -334 -1671 -332 -1667
rect -282 -1671 -280 -1667
rect -230 -1685 -228 -1676
rect -178 -1685 -176 -1676
rect 1262 -1657 1265 -1648
rect 1264 -1661 1265 -1657
rect 1262 -1676 1265 -1661
rect 1275 -1668 1278 -1648
rect 1339 -1667 1341 -1653
rect 1277 -1672 1278 -1668
rect 1275 -1676 1278 -1672
rect 1396 -1672 1398 -1669
rect 1406 -1672 1408 -1669
rect 1339 -1676 1341 -1673
rect -230 -1708 -228 -1705
rect -178 -1708 -176 -1705
rect -334 -1720 -332 -1711
rect -282 -1720 -280 -1711
rect -130 -1715 -128 -1695
rect -98 -1715 -96 -1695
rect 1262 -1697 1265 -1692
rect 1275 -1697 1278 -1692
rect 1437 -1685 1439 -1682
rect 1615 -1685 1617 -1682
rect 1625 -1685 1627 -1682
rect -334 -1732 -332 -1724
rect -282 -1732 -280 -1724
rect -230 -1732 -228 -1724
rect -178 -1732 -176 -1724
rect 1252 -1717 1255 -1713
rect 1265 -1717 1268 -1713
rect 1396 -1717 1398 -1696
rect 1406 -1717 1408 -1696
rect 1437 -1711 1439 -1697
rect 1656 -1698 1658 -1695
rect -130 -1739 -128 -1735
rect -98 -1739 -96 -1735
rect 1437 -1720 1439 -1717
rect 1396 -1726 1398 -1723
rect 1406 -1726 1408 -1723
rect 1329 -1730 1331 -1727
rect 1615 -1730 1617 -1709
rect 1625 -1730 1627 -1709
rect 1656 -1724 1658 -1710
rect 1252 -1746 1255 -1737
rect 1254 -1750 1255 -1746
rect -334 -1756 -332 -1752
rect -282 -1756 -280 -1752
rect -230 -1756 -228 -1752
rect -178 -1756 -176 -1752
rect 1252 -1765 1255 -1750
rect 1265 -1757 1268 -1737
rect 1656 -1733 1658 -1730
rect 1615 -1739 1617 -1736
rect 1625 -1739 1627 -1736
rect 1329 -1756 1331 -1742
rect 1267 -1761 1268 -1757
rect 1265 -1765 1268 -1761
rect 1329 -1765 1331 -1762
rect 1252 -1786 1255 -1781
rect 1265 -1786 1268 -1781
rect -334 -1832 -332 -1828
rect -282 -1832 -280 -1828
rect -230 -1832 -228 -1828
rect -178 -1832 -176 -1828
rect -334 -1881 -332 -1872
rect -282 -1881 -280 -1872
rect -230 -1881 -228 -1872
rect -178 -1881 -176 -1872
rect -130 -1878 -128 -1874
rect -98 -1878 -96 -1874
rect -334 -1894 -332 -1890
rect -282 -1894 -280 -1890
rect -230 -1908 -228 -1899
rect -178 -1908 -176 -1899
rect -230 -1931 -228 -1928
rect -178 -1931 -176 -1928
rect -334 -1943 -332 -1934
rect -282 -1943 -280 -1934
rect -130 -1938 -128 -1918
rect -98 -1938 -96 -1918
rect -334 -1955 -332 -1947
rect -282 -1955 -280 -1947
rect -230 -1955 -228 -1947
rect -178 -1955 -176 -1947
rect -130 -1962 -128 -1958
rect -98 -1962 -96 -1958
rect -334 -1979 -332 -1975
rect -282 -1979 -280 -1975
rect -230 -1979 -228 -1975
rect -178 -1979 -176 -1975
<< polycontact >>
rect -326 -315 -321 -310
rect -274 -315 -269 -310
rect -222 -315 -217 -310
rect -170 -315 -165 -310
rect -222 -338 -217 -333
rect -170 -338 -165 -333
rect 1581 -329 1586 -324
rect 1633 -329 1638 -324
rect 1685 -329 1690 -324
rect 1737 -329 1742 -324
rect -326 -377 -321 -372
rect -274 -377 -269 -372
rect -122 -369 -117 -364
rect -90 -369 -85 -364
rect -326 -386 -321 -381
rect -274 -386 -269 -381
rect -222 -386 -217 -381
rect -170 -386 -165 -381
rect 1685 -352 1690 -347
rect 1737 -352 1742 -347
rect 1581 -391 1586 -386
rect 1633 -391 1638 -386
rect 1785 -383 1790 -378
rect 1817 -383 1822 -378
rect 1581 -400 1586 -395
rect 1633 -400 1638 -395
rect 1685 -400 1690 -395
rect 1737 -400 1742 -395
rect 151 -480 155 -476
rect 182 -480 186 -476
rect 151 -530 155 -526
rect 192 -500 196 -496
rect -329 -542 -324 -537
rect -277 -542 -272 -537
rect -225 -542 -220 -537
rect -173 -542 -168 -537
rect -225 -565 -220 -560
rect -173 -565 -168 -560
rect 182 -553 186 -549
rect 202 -561 206 -557
rect 964 -550 968 -546
rect 995 -550 999 -546
rect -329 -604 -324 -599
rect -277 -604 -272 -599
rect -125 -596 -120 -591
rect -93 -596 -88 -591
rect -329 -613 -324 -608
rect -277 -613 -272 -608
rect -225 -613 -220 -608
rect -173 -613 -168 -608
rect 152 -601 156 -597
rect 183 -601 187 -597
rect 152 -651 156 -647
rect 193 -621 197 -617
rect 964 -600 968 -596
rect 1005 -570 1009 -566
rect 1573 -571 1578 -566
rect 1625 -571 1630 -566
rect 1677 -571 1682 -566
rect 1729 -571 1734 -566
rect 995 -623 999 -619
rect 183 -674 187 -670
rect 203 -682 207 -678
rect 637 -661 641 -657
rect 1015 -631 1019 -627
rect 1677 -594 1682 -589
rect 1729 -594 1734 -589
rect 1573 -633 1578 -628
rect 1625 -633 1630 -628
rect 1777 -625 1782 -620
rect 1809 -625 1814 -620
rect 1573 -642 1578 -637
rect 716 -664 720 -660
rect 649 -672 654 -668
rect 785 -671 789 -667
rect 795 -664 799 -660
rect 1625 -642 1630 -637
rect 1677 -642 1682 -637
rect 1729 -642 1734 -637
rect 826 -665 830 -661
rect 974 -674 978 -670
rect 1005 -674 1009 -670
rect 152 -722 156 -718
rect 183 -722 187 -718
rect -332 -771 -327 -766
rect -280 -771 -275 -766
rect -228 -771 -223 -766
rect -176 -771 -171 -766
rect -228 -794 -223 -789
rect -176 -794 -171 -789
rect 152 -772 156 -768
rect 193 -742 197 -738
rect 974 -724 978 -720
rect 1015 -694 1019 -690
rect 499 -754 504 -748
rect 511 -761 515 -757
rect 1005 -747 1009 -743
rect 555 -754 561 -749
rect 519 -768 523 -764
rect 183 -795 187 -791
rect 203 -803 207 -799
rect 1025 -755 1029 -751
rect 608 -791 612 -787
rect 618 -784 622 -780
rect 649 -785 653 -781
rect -332 -833 -327 -828
rect -280 -833 -275 -828
rect -128 -825 -123 -820
rect -96 -825 -91 -820
rect -332 -842 -327 -837
rect -280 -842 -275 -837
rect -228 -842 -223 -837
rect -176 -842 -171 -837
rect 152 -842 156 -838
rect 183 -842 187 -838
rect 152 -892 156 -888
rect 193 -862 197 -858
rect 878 -828 882 -824
rect 909 -828 913 -824
rect 498 -852 502 -848
rect 572 -855 576 -851
rect 510 -863 515 -859
rect 647 -899 651 -895
rect 183 -915 187 -911
rect 203 -923 207 -919
rect 657 -892 661 -888
rect 878 -878 882 -874
rect 919 -848 923 -844
rect 1574 -807 1579 -802
rect 1626 -807 1631 -802
rect 1678 -807 1683 -802
rect 1730 -807 1735 -802
rect 1678 -830 1683 -825
rect 1730 -830 1735 -825
rect 1574 -869 1579 -864
rect 1626 -869 1631 -864
rect 1778 -861 1783 -856
rect 1810 -861 1815 -856
rect 1574 -878 1579 -873
rect 1626 -878 1631 -873
rect 1678 -878 1683 -873
rect 1730 -878 1735 -873
rect 688 -893 692 -889
rect 909 -901 913 -897
rect 929 -909 933 -905
rect -332 -987 -327 -982
rect -280 -987 -275 -982
rect -228 -987 -223 -982
rect -176 -987 -171 -982
rect -228 -1010 -223 -1005
rect -176 -1010 -171 -1005
rect 856 -1022 860 -1018
rect -332 -1049 -327 -1044
rect -280 -1049 -275 -1044
rect -128 -1041 -123 -1036
rect -96 -1041 -91 -1036
rect 931 -1025 935 -1021
rect 868 -1033 873 -1029
rect -332 -1058 -327 -1053
rect -280 -1058 -275 -1053
rect -228 -1058 -223 -1053
rect -176 -1058 -171 -1053
rect 1574 -1040 1579 -1035
rect 1626 -1040 1631 -1035
rect 1678 -1040 1683 -1035
rect 1730 -1040 1735 -1035
rect 175 -1095 179 -1091
rect 250 -1098 254 -1094
rect 1007 -1094 1011 -1090
rect 187 -1106 192 -1102
rect 1017 -1087 1021 -1083
rect 1048 -1088 1052 -1084
rect 860 -1129 864 -1125
rect 1322 -1114 1326 -1110
rect 1353 -1114 1357 -1110
rect 935 -1132 939 -1128
rect 872 -1140 877 -1136
rect 176 -1182 180 -1178
rect -333 -1202 -328 -1197
rect -281 -1202 -276 -1197
rect -229 -1202 -224 -1197
rect -177 -1202 -172 -1197
rect 1095 -1173 1099 -1169
rect 250 -1185 254 -1181
rect 1105 -1166 1109 -1162
rect 1136 -1167 1140 -1163
rect 1322 -1164 1326 -1160
rect 1363 -1134 1367 -1130
rect 1678 -1063 1683 -1058
rect 1730 -1063 1735 -1058
rect 1574 -1102 1579 -1097
rect 1626 -1102 1631 -1097
rect 1778 -1094 1783 -1089
rect 1810 -1094 1815 -1089
rect 1574 -1111 1579 -1106
rect 1626 -1111 1631 -1106
rect 1678 -1111 1683 -1106
rect 1730 -1111 1735 -1106
rect 1353 -1187 1357 -1183
rect 188 -1193 193 -1189
rect 1373 -1195 1377 -1191
rect -229 -1225 -224 -1220
rect -177 -1225 -172 -1220
rect -333 -1264 -328 -1259
rect -281 -1264 -276 -1259
rect -129 -1256 -124 -1251
rect -97 -1256 -92 -1251
rect 860 -1238 864 -1234
rect -333 -1273 -328 -1268
rect -281 -1273 -276 -1268
rect -229 -1273 -224 -1268
rect -177 -1273 -172 -1268
rect 178 -1270 182 -1266
rect 935 -1241 939 -1237
rect 872 -1249 877 -1245
rect 253 -1273 257 -1269
rect 1007 -1263 1011 -1259
rect 1017 -1256 1021 -1252
rect 1048 -1257 1052 -1253
rect 1569 -1266 1574 -1261
rect 1621 -1266 1626 -1261
rect 1673 -1266 1678 -1261
rect 1725 -1266 1730 -1261
rect 190 -1281 195 -1277
rect 1673 -1289 1678 -1284
rect 1725 -1289 1730 -1284
rect 1569 -1328 1574 -1323
rect 1621 -1328 1626 -1323
rect 1773 -1320 1778 -1315
rect 1805 -1320 1810 -1315
rect 178 -1356 182 -1352
rect 1569 -1337 1574 -1332
rect 1621 -1337 1626 -1332
rect 1673 -1337 1678 -1332
rect 1725 -1337 1730 -1332
rect 254 -1359 258 -1355
rect 190 -1367 195 -1363
rect -341 -1432 -336 -1427
rect -289 -1432 -284 -1427
rect -237 -1432 -232 -1427
rect -185 -1432 -180 -1427
rect -237 -1455 -232 -1450
rect -185 -1455 -180 -1450
rect 1260 -1453 1264 -1449
rect 1335 -1456 1339 -1452
rect 1272 -1464 1277 -1460
rect -341 -1494 -336 -1489
rect -289 -1494 -284 -1489
rect -137 -1486 -132 -1481
rect -105 -1486 -100 -1481
rect -341 -1503 -336 -1498
rect -289 -1503 -284 -1498
rect -237 -1503 -232 -1498
rect -185 -1503 -180 -1498
rect 1395 -1512 1399 -1508
rect 1405 -1505 1409 -1501
rect 1436 -1506 1440 -1502
rect 1260 -1558 1264 -1554
rect 1335 -1561 1339 -1557
rect 1272 -1569 1277 -1565
rect 1508 -1625 1512 -1621
rect 1518 -1618 1522 -1614
rect 1549 -1619 1553 -1615
rect -339 -1658 -334 -1653
rect -287 -1658 -282 -1653
rect -235 -1658 -230 -1653
rect -183 -1658 -178 -1653
rect -235 -1681 -230 -1676
rect -183 -1681 -178 -1676
rect 1260 -1661 1264 -1657
rect 1335 -1664 1339 -1660
rect 1272 -1672 1277 -1668
rect -339 -1720 -334 -1715
rect -287 -1720 -282 -1715
rect -135 -1712 -130 -1707
rect -103 -1712 -98 -1707
rect -339 -1729 -334 -1724
rect -287 -1729 -282 -1724
rect -235 -1729 -230 -1724
rect -183 -1729 -178 -1724
rect 1392 -1714 1396 -1710
rect 1402 -1707 1406 -1703
rect 1433 -1708 1437 -1704
rect 1611 -1727 1615 -1723
rect 1621 -1720 1625 -1716
rect 1652 -1721 1656 -1717
rect 1250 -1750 1254 -1746
rect 1325 -1753 1329 -1749
rect 1262 -1761 1267 -1757
rect -339 -1881 -334 -1876
rect -287 -1881 -282 -1876
rect -235 -1881 -230 -1876
rect -183 -1881 -178 -1876
rect -235 -1904 -230 -1899
rect -183 -1904 -178 -1899
rect -339 -1943 -334 -1938
rect -287 -1943 -282 -1938
rect -135 -1935 -130 -1930
rect -103 -1935 -98 -1930
rect -339 -1952 -334 -1947
rect -287 -1952 -282 -1947
rect -235 -1952 -230 -1947
rect -183 -1952 -178 -1947
<< metal1 >>
rect -336 -254 -148 -251
rect -336 -258 -333 -254
rect -329 -258 -311 -254
rect -307 -258 -281 -254
rect -277 -258 -259 -254
rect -255 -258 -229 -254
rect -225 -258 -207 -254
rect -203 -258 -177 -254
rect -173 -258 -155 -254
rect -151 -258 -148 -254
rect -336 -260 -148 -258
rect -326 -266 -322 -260
rect -274 -266 -270 -260
rect -222 -266 -218 -260
rect -170 -266 -166 -260
rect 1571 -268 1759 -265
rect 1571 -272 1574 -268
rect 1578 -272 1596 -268
rect 1600 -272 1626 -268
rect 1630 -272 1648 -268
rect 1652 -272 1678 -268
rect 1682 -272 1700 -268
rect 1704 -272 1730 -268
rect 1734 -272 1752 -268
rect 1756 -272 1759 -268
rect 1571 -274 1759 -272
rect 1581 -280 1585 -274
rect 1633 -280 1637 -274
rect 1685 -280 1689 -274
rect 1737 -280 1741 -274
rect -132 -300 -68 -297
rect -132 -304 -129 -300
rect -125 -304 -107 -300
rect -103 -304 -97 -300
rect -93 -304 -75 -300
rect -71 -304 -68 -300
rect -132 -306 -68 -304
rect -349 -315 -326 -310
rect -349 -344 -344 -315
rect -318 -319 -314 -306
rect -362 -349 -344 -344
rect -349 -381 -344 -349
rect -326 -323 -314 -319
rect -296 -315 -274 -310
rect -326 -328 -322 -323
rect -331 -377 -326 -372
rect -318 -381 -314 -368
rect -296 -381 -291 -315
rect -266 -319 -262 -306
rect -214 -310 -210 -306
rect -162 -310 -158 -306
rect -274 -323 -262 -319
rect -244 -315 -222 -310
rect -214 -315 -170 -310
rect -162 -315 -142 -310
rect -274 -328 -270 -323
rect -279 -377 -274 -372
rect -266 -381 -262 -368
rect -244 -381 -239 -315
rect -225 -338 -222 -333
rect -214 -342 -210 -315
rect -222 -373 -218 -362
rect -222 -377 -210 -373
rect -349 -386 -326 -381
rect -318 -386 -274 -381
rect -266 -386 -222 -381
rect -318 -389 -314 -386
rect -266 -389 -262 -386
rect -214 -389 -210 -377
rect -192 -381 -187 -315
rect -173 -338 -170 -333
rect -162 -342 -158 -315
rect -170 -373 -166 -362
rect -147 -364 -142 -315
rect -122 -312 -118 -306
rect -90 -312 -86 -306
rect 1775 -314 1839 -311
rect 1775 -318 1778 -314
rect 1782 -318 1800 -314
rect 1804 -318 1810 -314
rect 1814 -318 1832 -314
rect 1836 -318 1839 -314
rect 1775 -320 1839 -318
rect -114 -364 -110 -352
rect -82 -364 -78 -352
rect 1558 -329 1581 -324
rect 1558 -358 1563 -329
rect 1589 -333 1593 -320
rect 1545 -363 1563 -358
rect -147 -369 -122 -364
rect -114 -369 -90 -364
rect -82 -369 -48 -364
rect -114 -372 -110 -369
rect -82 -372 -78 -369
rect -170 -377 -158 -373
rect -192 -386 -170 -381
rect -162 -389 -158 -377
rect -122 -399 -118 -392
rect -90 -399 -86 -392
rect 1558 -395 1563 -363
rect 1581 -337 1593 -333
rect 1611 -329 1633 -324
rect 1581 -342 1585 -337
rect 1576 -391 1581 -386
rect 1589 -395 1593 -382
rect 1611 -395 1616 -329
rect 1641 -333 1645 -320
rect 1693 -324 1697 -320
rect 1745 -324 1749 -320
rect 1633 -337 1645 -333
rect 1663 -329 1685 -324
rect 1693 -329 1737 -324
rect 1745 -329 1765 -324
rect 1633 -342 1637 -337
rect 1628 -391 1633 -386
rect 1641 -395 1645 -382
rect 1663 -395 1668 -329
rect 1682 -352 1685 -347
rect 1693 -356 1697 -329
rect 1685 -387 1689 -376
rect 1685 -391 1697 -387
rect -132 -401 -68 -399
rect 1558 -400 1581 -395
rect 1589 -400 1633 -395
rect 1641 -400 1685 -395
rect -132 -405 -130 -401
rect -126 -405 -106 -401
rect -102 -405 -98 -401
rect -94 -405 -74 -401
rect -70 -405 -68 -401
rect 1589 -403 1593 -400
rect 1641 -403 1645 -400
rect 1693 -403 1697 -391
rect 1715 -395 1720 -329
rect 1734 -352 1737 -347
rect 1745 -356 1749 -329
rect 1737 -387 1741 -376
rect 1760 -378 1765 -329
rect 1785 -326 1789 -320
rect 1817 -326 1821 -320
rect 1793 -378 1797 -366
rect 1825 -378 1829 -366
rect 1760 -383 1785 -378
rect 1793 -383 1817 -378
rect 1825 -383 1859 -378
rect 1793 -386 1797 -383
rect 1825 -386 1829 -383
rect 1737 -391 1749 -387
rect 1715 -400 1737 -395
rect 1745 -403 1749 -391
rect -132 -407 -68 -405
rect -326 -417 -322 -409
rect -274 -417 -270 -409
rect -222 -417 -218 -409
rect -170 -417 -166 -409
rect -336 -418 -148 -417
rect -336 -422 -309 -418
rect -305 -422 -257 -418
rect -253 -422 -205 -418
rect -201 -422 -153 -418
rect -149 -422 -148 -418
rect -336 -423 -148 -422
rect 1785 -413 1789 -406
rect 1817 -413 1821 -406
rect 1775 -415 1839 -413
rect 1775 -419 1777 -415
rect 1781 -419 1801 -415
rect 1805 -419 1809 -415
rect 1813 -419 1833 -415
rect 1837 -419 1839 -415
rect 1775 -421 1839 -419
rect 1581 -431 1585 -423
rect 1633 -431 1637 -423
rect 1685 -431 1689 -423
rect 1737 -431 1741 -423
rect -343 -436 -336 -431
rect -331 -436 -284 -431
rect -279 -436 -230 -431
rect -225 -436 -178 -431
rect 1571 -432 1759 -431
rect 1571 -436 1598 -432
rect 1602 -436 1650 -432
rect 1654 -436 1702 -432
rect 1706 -436 1754 -432
rect 1758 -436 1759 -432
rect 1571 -437 1759 -436
rect 1564 -450 1571 -445
rect 1576 -450 1623 -445
rect 1628 -450 1677 -445
rect 1682 -450 1729 -445
rect 121 -455 230 -451
rect -339 -481 -151 -478
rect 14 -480 125 -476
rect -339 -485 -336 -481
rect -332 -485 -314 -481
rect -310 -485 -284 -481
rect -280 -485 -262 -481
rect -258 -485 -232 -481
rect -228 -485 -210 -481
rect -206 -485 -180 -481
rect -176 -485 -158 -481
rect -154 -485 -151 -481
rect -339 -487 -151 -485
rect -329 -493 -325 -487
rect -277 -493 -273 -487
rect -225 -493 -221 -487
rect -173 -493 -169 -487
rect 135 -501 139 -455
rect 150 -461 154 -455
rect 180 -461 184 -455
rect 220 -461 224 -455
rect 158 -476 162 -469
rect 147 -480 151 -476
rect 158 -480 182 -476
rect 158 -483 162 -480
rect 150 -491 154 -487
rect 144 -495 177 -491
rect 135 -505 168 -501
rect 150 -511 154 -505
rect -135 -527 -71 -524
rect 158 -526 162 -519
rect -135 -531 -132 -527
rect -128 -531 -110 -527
rect -106 -531 -100 -527
rect -96 -531 -78 -527
rect -74 -531 -71 -527
rect 13 -530 134 -526
rect 139 -530 151 -526
rect 158 -530 165 -526
rect -135 -533 -71 -531
rect 158 -533 162 -530
rect -352 -542 -329 -537
rect -352 -571 -347 -542
rect -321 -546 -317 -533
rect -365 -576 -347 -571
rect -352 -608 -347 -576
rect -329 -550 -317 -546
rect -299 -542 -277 -537
rect -329 -555 -325 -550
rect -334 -604 -329 -599
rect -321 -608 -317 -595
rect -299 -608 -294 -542
rect -269 -546 -265 -533
rect -217 -537 -213 -533
rect -165 -537 -161 -533
rect -277 -550 -265 -546
rect -247 -542 -225 -537
rect -217 -542 -173 -537
rect -165 -542 -145 -537
rect -277 -555 -273 -550
rect -282 -604 -277 -599
rect -269 -608 -265 -595
rect -247 -608 -242 -542
rect -228 -565 -225 -560
rect -217 -569 -213 -542
rect -225 -600 -221 -589
rect -225 -604 -213 -600
rect -352 -613 -329 -608
rect -321 -613 -277 -608
rect -269 -613 -225 -608
rect -321 -616 -317 -613
rect -269 -616 -265 -613
rect -217 -616 -213 -604
rect -195 -608 -190 -542
rect -176 -565 -173 -560
rect -165 -569 -161 -542
rect -173 -600 -169 -589
rect -150 -591 -145 -542
rect -125 -539 -121 -533
rect -93 -539 -89 -533
rect 150 -541 154 -537
rect 173 -541 177 -495
rect 185 -500 192 -496
rect 200 -502 204 -469
rect 200 -506 908 -502
rect 200 -533 204 -506
rect 180 -541 184 -537
rect 220 -541 224 -537
rect 121 -545 230 -541
rect 140 -553 182 -549
rect 171 -561 202 -557
rect 122 -576 231 -572
rect -117 -591 -113 -579
rect -85 -591 -81 -579
rect -150 -596 -125 -591
rect -117 -596 -93 -591
rect -85 -596 -51 -591
rect -117 -599 -113 -596
rect -85 -599 -81 -596
rect -173 -604 -161 -600
rect -195 -613 -173 -608
rect -165 -616 -161 -604
rect 15 -601 126 -597
rect -125 -626 -121 -619
rect -93 -626 -89 -619
rect 136 -622 140 -576
rect 151 -582 155 -576
rect 181 -582 185 -576
rect 221 -582 225 -576
rect 159 -597 163 -590
rect 148 -601 152 -597
rect 159 -601 183 -597
rect 159 -604 163 -601
rect 151 -612 155 -608
rect 145 -616 178 -612
rect 136 -626 169 -622
rect -135 -628 -71 -626
rect -135 -632 -133 -628
rect -129 -632 -109 -628
rect -105 -632 -101 -628
rect -97 -632 -77 -628
rect -73 -632 -71 -628
rect -135 -634 -71 -632
rect 151 -632 155 -626
rect -329 -644 -325 -636
rect -277 -644 -273 -636
rect -225 -644 -221 -636
rect -173 -644 -169 -636
rect -339 -645 -151 -644
rect -339 -649 -312 -645
rect -308 -649 -260 -645
rect -256 -649 -208 -645
rect -204 -649 -156 -645
rect -152 -649 -151 -645
rect 159 -647 163 -640
rect -339 -650 -151 -649
rect 14 -651 135 -647
rect 140 -651 152 -647
rect 159 -651 166 -647
rect 159 -654 163 -651
rect -346 -663 -339 -658
rect -334 -663 -287 -658
rect -282 -663 -233 -658
rect -228 -663 -181 -658
rect 151 -662 155 -658
rect 174 -662 178 -616
rect 186 -621 193 -617
rect 201 -623 205 -590
rect 374 -623 378 -616
rect 201 -627 441 -623
rect 201 -654 205 -627
rect 181 -662 185 -658
rect 221 -662 225 -658
rect 122 -666 231 -662
rect 141 -674 183 -670
rect 172 -682 203 -678
rect 122 -697 231 -693
rect -342 -710 -154 -707
rect -342 -714 -339 -710
rect -335 -714 -317 -710
rect -313 -714 -287 -710
rect -283 -714 -265 -710
rect -261 -714 -235 -710
rect -231 -714 -213 -710
rect -209 -714 -183 -710
rect -179 -714 -161 -710
rect -157 -714 -154 -710
rect -342 -716 -154 -714
rect -332 -722 -328 -716
rect -280 -722 -276 -716
rect -228 -722 -224 -716
rect -176 -722 -172 -716
rect 15 -722 126 -718
rect 136 -743 140 -697
rect 151 -703 155 -697
rect 181 -703 185 -697
rect 221 -703 225 -697
rect 159 -718 163 -711
rect 148 -722 152 -718
rect 159 -722 183 -718
rect 159 -725 163 -722
rect 151 -733 155 -729
rect 145 -737 178 -733
rect 136 -747 169 -743
rect 151 -753 155 -747
rect -138 -756 -74 -753
rect -138 -760 -135 -756
rect -131 -760 -113 -756
rect -109 -760 -103 -756
rect -99 -760 -81 -756
rect -77 -760 -74 -756
rect -138 -762 -74 -760
rect -355 -771 -332 -766
rect -355 -800 -350 -771
rect -324 -775 -320 -762
rect -368 -805 -350 -800
rect -355 -837 -350 -805
rect -332 -779 -320 -775
rect -302 -771 -280 -766
rect -332 -784 -328 -779
rect -337 -833 -332 -828
rect -324 -837 -320 -824
rect -302 -837 -297 -771
rect -272 -775 -268 -762
rect -220 -766 -216 -762
rect -168 -766 -164 -762
rect -280 -779 -268 -775
rect -250 -771 -228 -766
rect -220 -771 -176 -766
rect -168 -771 -148 -766
rect -280 -784 -276 -779
rect -285 -833 -280 -828
rect -272 -837 -268 -824
rect -250 -837 -245 -771
rect -231 -794 -228 -789
rect -220 -798 -216 -771
rect -228 -829 -224 -818
rect -228 -833 -216 -829
rect -355 -842 -332 -837
rect -324 -842 -280 -837
rect -272 -842 -228 -837
rect -324 -845 -320 -842
rect -272 -845 -268 -842
rect -220 -845 -216 -833
rect -198 -837 -193 -771
rect -179 -794 -176 -789
rect -168 -798 -164 -771
rect -176 -829 -172 -818
rect -153 -820 -148 -771
rect -128 -768 -124 -762
rect -96 -768 -92 -762
rect 159 -768 163 -761
rect 14 -772 135 -768
rect 140 -772 152 -768
rect 159 -772 166 -768
rect 159 -775 163 -772
rect 151 -783 155 -779
rect 174 -783 178 -737
rect 186 -742 193 -738
rect 201 -744 205 -711
rect 321 -744 325 -693
rect 201 -748 370 -744
rect 201 -775 205 -748
rect 181 -783 185 -779
rect 221 -783 225 -779
rect 122 -787 231 -783
rect 141 -795 183 -791
rect 172 -803 203 -799
rect -120 -820 -116 -808
rect -88 -820 -84 -808
rect 122 -817 231 -813
rect -153 -825 -128 -820
rect -120 -825 -96 -820
rect -88 -825 -54 -820
rect -120 -828 -116 -825
rect -88 -828 -84 -825
rect -176 -833 -164 -829
rect -198 -842 -176 -837
rect -168 -845 -164 -833
rect 15 -842 126 -838
rect -128 -855 -124 -848
rect -96 -855 -92 -848
rect -138 -857 -74 -855
rect -138 -861 -136 -857
rect -132 -861 -112 -857
rect -108 -861 -104 -857
rect -100 -861 -80 -857
rect -76 -861 -74 -857
rect -138 -863 -74 -861
rect 136 -863 140 -817
rect 151 -823 155 -817
rect 181 -823 185 -817
rect 221 -823 225 -817
rect 159 -838 163 -831
rect 148 -842 152 -838
rect 159 -842 183 -838
rect 159 -845 163 -842
rect 151 -853 155 -849
rect 145 -857 178 -853
rect -332 -873 -328 -865
rect -280 -873 -276 -865
rect -228 -873 -224 -865
rect -176 -873 -172 -865
rect 136 -867 169 -863
rect 151 -873 155 -867
rect -342 -874 -154 -873
rect -342 -878 -315 -874
rect -311 -878 -263 -874
rect -259 -878 -211 -874
rect -207 -878 -159 -874
rect -155 -878 -154 -874
rect -342 -879 -154 -878
rect -349 -892 -342 -887
rect -337 -892 -290 -887
rect -285 -892 -236 -887
rect -231 -892 -184 -887
rect 159 -888 163 -881
rect 14 -892 135 -888
rect 140 -892 152 -888
rect 159 -892 166 -888
rect 159 -895 163 -892
rect 151 -903 155 -899
rect 174 -903 178 -857
rect 186 -862 193 -858
rect 201 -864 205 -831
rect 201 -868 325 -864
rect 201 -895 205 -868
rect 181 -903 185 -899
rect 221 -903 225 -899
rect 122 -907 231 -903
rect 141 -915 183 -911
rect 172 -923 203 -919
rect -342 -926 -154 -923
rect -342 -930 -339 -926
rect -335 -930 -317 -926
rect -313 -930 -287 -926
rect -283 -930 -265 -926
rect -261 -930 -235 -926
rect -231 -930 -213 -926
rect -209 -930 -183 -926
rect -179 -930 -161 -926
rect -157 -930 -154 -926
rect -342 -932 -154 -930
rect -332 -938 -328 -932
rect -280 -938 -276 -932
rect -228 -938 -224 -932
rect -176 -938 -172 -932
rect -138 -972 -74 -969
rect -138 -976 -135 -972
rect -131 -976 -113 -972
rect -109 -976 -103 -972
rect -99 -976 -81 -972
rect -77 -976 -74 -972
rect -138 -978 -74 -976
rect -355 -987 -332 -982
rect -355 -1016 -350 -987
rect -324 -991 -320 -978
rect -368 -1021 -350 -1016
rect -355 -1053 -350 -1021
rect -332 -995 -320 -991
rect -302 -987 -280 -982
rect -332 -1000 -328 -995
rect -337 -1049 -332 -1044
rect -324 -1053 -320 -1040
rect -302 -1053 -297 -987
rect -272 -991 -268 -978
rect -220 -982 -216 -978
rect -168 -982 -164 -978
rect -280 -995 -268 -991
rect -250 -987 -228 -982
rect -220 -987 -176 -982
rect -168 -987 -148 -982
rect -280 -1000 -276 -995
rect -285 -1049 -280 -1044
rect -272 -1053 -268 -1040
rect -250 -1053 -245 -987
rect -231 -1010 -228 -1005
rect -220 -1014 -216 -987
rect -228 -1045 -224 -1034
rect -228 -1049 -216 -1045
rect -355 -1058 -332 -1053
rect -324 -1058 -280 -1053
rect -272 -1058 -228 -1053
rect -324 -1061 -320 -1058
rect -272 -1061 -268 -1058
rect -220 -1061 -216 -1049
rect -198 -1053 -193 -987
rect -179 -1010 -176 -1005
rect -168 -1014 -164 -987
rect -176 -1045 -172 -1034
rect -153 -1036 -148 -987
rect -128 -984 -124 -978
rect -96 -984 -92 -978
rect -120 -1036 -116 -1024
rect -88 -1036 -84 -1024
rect 321 -993 325 -868
rect 321 -997 332 -993
rect -153 -1041 -128 -1036
rect -120 -1041 -96 -1036
rect -88 -1041 -54 -1036
rect -120 -1044 -116 -1041
rect -88 -1044 -84 -1041
rect -176 -1049 -164 -1045
rect -198 -1058 -176 -1053
rect -168 -1061 -164 -1049
rect 171 -1054 199 -1050
rect 171 -1062 175 -1054
rect 195 -1062 199 -1054
rect -128 -1071 -124 -1064
rect -96 -1071 -92 -1064
rect -138 -1073 -74 -1071
rect -138 -1077 -136 -1073
rect -132 -1077 -112 -1073
rect -108 -1077 -104 -1073
rect -100 -1077 -80 -1073
rect -76 -1077 -74 -1073
rect -138 -1079 -74 -1077
rect -332 -1089 -328 -1081
rect -280 -1089 -276 -1081
rect -228 -1089 -224 -1081
rect -176 -1089 -172 -1081
rect -342 -1090 -154 -1089
rect -342 -1094 -315 -1090
rect -311 -1094 -263 -1090
rect -259 -1094 -211 -1090
rect -207 -1094 -159 -1090
rect -155 -1094 -154 -1090
rect -342 -1095 -154 -1094
rect 115 -1095 175 -1091
rect 183 -1095 187 -1067
rect 243 -1069 267 -1066
rect 321 -1069 325 -997
rect 366 -1021 370 -748
rect 437 -764 441 -627
rect 450 -757 454 -506
rect 571 -550 575 -506
rect 904 -546 908 -506
rect 1563 -510 1751 -507
rect 1563 -514 1566 -510
rect 1570 -514 1588 -510
rect 1592 -514 1618 -510
rect 1622 -514 1640 -510
rect 1644 -514 1670 -510
rect 1674 -514 1692 -510
rect 1696 -514 1722 -510
rect 1726 -514 1744 -510
rect 1748 -514 1751 -510
rect 1563 -516 1751 -514
rect 934 -525 1043 -521
rect 1573 -522 1577 -516
rect 1625 -522 1629 -516
rect 1677 -522 1681 -516
rect 1729 -522 1733 -516
rect 904 -550 938 -546
rect 537 -562 563 -557
rect 537 -668 542 -562
rect 571 -654 575 -564
rect 885 -562 898 -558
rect 894 -596 898 -562
rect 948 -571 952 -525
rect 963 -531 967 -525
rect 993 -531 997 -525
rect 1033 -531 1037 -525
rect 971 -546 975 -539
rect 960 -550 964 -546
rect 971 -550 995 -546
rect 971 -553 975 -550
rect 963 -561 967 -557
rect 957 -565 990 -561
rect 948 -575 981 -571
rect 963 -581 967 -575
rect 971 -596 975 -589
rect 894 -600 947 -596
rect 952 -600 964 -596
rect 971 -600 978 -596
rect 971 -603 975 -600
rect 963 -611 967 -607
rect 986 -611 990 -565
rect 998 -570 1005 -566
rect 1013 -572 1017 -539
rect 1767 -556 1831 -553
rect 1767 -560 1770 -556
rect 1774 -560 1792 -556
rect 1796 -560 1802 -556
rect 1806 -560 1824 -556
rect 1828 -560 1831 -556
rect 1767 -562 1831 -560
rect 1550 -571 1573 -566
rect 1013 -576 1111 -572
rect 1013 -603 1017 -576
rect 1550 -600 1555 -571
rect 1581 -575 1585 -562
rect 1537 -605 1555 -600
rect 993 -611 997 -607
rect 1033 -611 1037 -607
rect 934 -615 1043 -611
rect 633 -620 661 -616
rect 633 -628 637 -620
rect 657 -628 661 -620
rect 778 -623 812 -620
rect 953 -623 995 -619
rect 784 -629 787 -623
rect 570 -657 618 -654
rect 570 -661 637 -657
rect 645 -661 649 -633
rect 709 -635 733 -632
rect 715 -641 718 -635
rect 984 -631 1015 -627
rect 819 -636 843 -633
rect 655 -661 710 -660
rect 645 -664 716 -661
rect 724 -661 727 -653
rect 730 -661 765 -660
rect 724 -664 795 -661
rect 803 -662 806 -653
rect 825 -642 828 -636
rect 1550 -637 1555 -605
rect 1573 -579 1585 -575
rect 1603 -571 1625 -566
rect 1573 -584 1577 -579
rect 1568 -633 1573 -628
rect 1581 -637 1585 -624
rect 1603 -637 1608 -571
rect 1633 -575 1637 -562
rect 1685 -566 1689 -562
rect 1737 -566 1741 -562
rect 1625 -579 1637 -575
rect 1655 -571 1677 -566
rect 1685 -571 1729 -566
rect 1737 -571 1757 -566
rect 1625 -584 1629 -579
rect 1620 -633 1625 -628
rect 1633 -637 1637 -624
rect 1655 -637 1660 -571
rect 1674 -594 1677 -589
rect 1685 -598 1689 -571
rect 1677 -629 1681 -618
rect 1677 -633 1689 -629
rect 1550 -642 1573 -637
rect 1581 -642 1625 -637
rect 1633 -642 1677 -637
rect 1581 -645 1585 -642
rect 1633 -645 1637 -642
rect 1685 -645 1689 -633
rect 1707 -637 1712 -571
rect 1726 -594 1729 -589
rect 1737 -598 1741 -571
rect 1729 -629 1733 -618
rect 1752 -620 1757 -571
rect 1777 -568 1781 -562
rect 1809 -568 1813 -562
rect 1785 -620 1789 -608
rect 1817 -620 1821 -608
rect 1752 -625 1777 -620
rect 1785 -625 1809 -620
rect 1817 -625 1851 -620
rect 1785 -628 1789 -625
rect 1817 -628 1821 -625
rect 1729 -633 1741 -629
rect 1707 -642 1729 -637
rect 1737 -645 1741 -633
rect 944 -649 1053 -645
rect 645 -665 710 -664
rect 464 -672 649 -668
rect 654 -672 655 -668
rect 464 -673 655 -672
rect 464 -748 469 -673
rect 658 -676 661 -665
rect 724 -667 727 -664
rect 730 -665 755 -664
rect 803 -665 826 -662
rect 834 -662 837 -654
rect 843 -662 898 -661
rect 834 -665 898 -662
rect 759 -670 785 -667
rect 715 -677 718 -673
rect 709 -680 733 -677
rect 633 -696 637 -681
rect 495 -700 532 -699
rect 495 -704 497 -700
rect 501 -704 509 -700
rect 513 -704 518 -700
rect 522 -704 526 -700
rect 530 -704 532 -700
rect 495 -706 532 -704
rect 547 -706 577 -703
rect 496 -714 500 -706
rect 516 -714 520 -706
rect 547 -710 550 -706
rect 554 -710 558 -706
rect 562 -710 566 -706
rect 570 -710 577 -706
rect 547 -711 577 -710
rect 554 -717 559 -711
rect 582 -725 730 -722
rect 464 -753 499 -748
rect 498 -754 499 -753
rect 507 -750 511 -739
rect 527 -749 531 -739
rect 527 -750 555 -749
rect 507 -754 555 -750
rect 564 -750 569 -737
rect 582 -750 585 -725
rect 601 -743 635 -740
rect 607 -749 610 -743
rect 564 -753 594 -750
rect 450 -761 511 -757
rect 437 -768 519 -764
rect 437 -848 441 -768
rect 527 -771 531 -754
rect 564 -758 569 -753
rect 555 -774 559 -768
rect 546 -777 580 -774
rect 496 -789 501 -781
rect 546 -782 549 -777
rect 572 -782 580 -777
rect 546 -784 580 -782
rect 591 -781 594 -753
rect 642 -756 666 -753
rect 591 -784 618 -781
rect 626 -782 629 -773
rect 648 -762 651 -756
rect 626 -785 649 -782
rect 657 -782 660 -774
rect 657 -785 673 -782
rect 495 -790 532 -789
rect 495 -794 497 -790
rect 501 -794 505 -790
rect 509 -794 513 -790
rect 517 -794 521 -790
rect 525 -794 532 -790
rect 495 -796 532 -794
rect 595 -790 608 -787
rect 494 -811 522 -807
rect 494 -819 498 -811
rect 518 -819 522 -811
rect 437 -852 498 -848
rect 506 -852 510 -824
rect 565 -826 589 -823
rect 571 -832 574 -826
rect 516 -852 566 -851
rect 506 -855 572 -852
rect 580 -852 583 -844
rect 595 -851 598 -790
rect 626 -788 629 -785
rect 657 -788 660 -785
rect 617 -791 629 -788
rect 617 -794 620 -791
rect 648 -798 651 -794
rect 607 -806 610 -800
rect 626 -806 629 -800
rect 642 -801 666 -798
rect 601 -809 635 -806
rect 670 -827 673 -785
rect 586 -852 598 -851
rect 580 -855 598 -852
rect 506 -856 566 -855
rect 438 -863 510 -859
rect 515 -863 516 -859
rect 438 -864 516 -863
rect 249 -1075 252 -1069
rect 317 -1071 338 -1069
rect 193 -1095 244 -1094
rect 183 -1098 250 -1095
rect 258 -1095 261 -1087
rect 438 -1094 443 -864
rect 519 -867 522 -856
rect 580 -858 583 -855
rect 586 -856 598 -855
rect 613 -830 673 -827
rect 571 -868 574 -864
rect 565 -871 589 -868
rect 494 -887 498 -872
rect 592 -879 597 -856
rect 535 -884 597 -879
rect 535 -1047 540 -884
rect 613 -889 616 -830
rect 640 -851 674 -848
rect 646 -857 649 -851
rect 681 -864 705 -861
rect 613 -892 657 -889
rect 665 -890 668 -881
rect 687 -870 690 -864
rect 665 -893 688 -890
rect 696 -890 699 -882
rect 696 -893 723 -890
rect 553 -898 647 -895
rect 553 -1063 556 -898
rect 665 -896 668 -893
rect 696 -896 699 -893
rect 656 -899 668 -896
rect 656 -902 659 -899
rect 687 -906 690 -902
rect 646 -914 649 -908
rect 665 -914 668 -908
rect 681 -909 705 -906
rect 640 -917 674 -914
rect 551 -1074 558 -1063
rect 759 -1084 762 -670
rect 803 -668 806 -665
rect 834 -668 837 -665
rect 794 -671 806 -668
rect 794 -674 797 -671
rect 825 -678 828 -674
rect 784 -686 787 -680
rect 803 -686 806 -680
rect 819 -681 843 -678
rect 778 -689 812 -686
rect 894 -721 898 -665
rect 938 -674 948 -670
rect 958 -695 962 -649
rect 973 -655 977 -649
rect 1003 -655 1007 -649
rect 1043 -655 1047 -649
rect 981 -670 985 -663
rect 970 -674 974 -670
rect 981 -674 1005 -670
rect 981 -677 985 -674
rect 973 -685 977 -681
rect 967 -689 1000 -685
rect 958 -699 991 -695
rect 973 -705 977 -699
rect 981 -720 985 -713
rect 938 -721 957 -720
rect 894 -724 957 -721
rect 894 -725 941 -724
rect 962 -724 974 -720
rect 981 -724 988 -720
rect 981 -727 985 -724
rect 782 -853 793 -734
rect 973 -735 977 -731
rect 996 -735 1000 -689
rect 1008 -694 1015 -690
rect 1023 -696 1027 -663
rect 1777 -655 1781 -648
rect 1809 -655 1813 -648
rect 1767 -657 1831 -655
rect 1767 -661 1769 -657
rect 1773 -661 1793 -657
rect 1797 -661 1801 -657
rect 1805 -661 1825 -657
rect 1829 -661 1831 -657
rect 1767 -663 1831 -661
rect 1573 -673 1577 -665
rect 1625 -673 1629 -665
rect 1677 -673 1681 -665
rect 1729 -673 1733 -665
rect 1563 -674 1751 -673
rect 1563 -678 1590 -674
rect 1594 -678 1642 -674
rect 1646 -678 1694 -674
rect 1698 -678 1746 -674
rect 1750 -678 1751 -674
rect 1563 -679 1751 -678
rect 1556 -692 1563 -687
rect 1568 -692 1615 -687
rect 1620 -692 1669 -687
rect 1674 -692 1721 -687
rect 1023 -700 1087 -696
rect 1023 -727 1027 -700
rect 1003 -735 1007 -731
rect 1043 -735 1047 -731
rect 944 -739 1053 -735
rect 963 -747 1005 -743
rect 1564 -746 1752 -743
rect 1564 -750 1567 -746
rect 1571 -750 1589 -746
rect 1593 -750 1619 -746
rect 1623 -750 1641 -746
rect 1645 -750 1671 -746
rect 1675 -750 1693 -746
rect 1697 -750 1723 -746
rect 1727 -750 1745 -746
rect 1749 -750 1752 -746
rect 994 -755 1025 -751
rect 1564 -752 1752 -750
rect 1574 -758 1578 -752
rect 1626 -758 1630 -752
rect 1678 -758 1682 -752
rect 1730 -758 1734 -752
rect 1768 -792 1832 -789
rect 1768 -796 1771 -792
rect 1775 -796 1793 -792
rect 1797 -796 1803 -792
rect 1807 -796 1825 -792
rect 1829 -796 1832 -792
rect 1768 -798 1832 -796
rect 848 -803 957 -799
rect 839 -828 852 -824
rect 862 -849 866 -803
rect 877 -809 881 -803
rect 907 -809 911 -803
rect 947 -809 951 -803
rect 1551 -807 1574 -802
rect 885 -824 889 -817
rect 874 -828 878 -824
rect 885 -828 909 -824
rect 885 -831 889 -828
rect 877 -839 881 -835
rect 871 -843 904 -839
rect 862 -853 895 -849
rect 788 -1018 792 -853
rect 877 -859 881 -853
rect 885 -874 889 -867
rect 838 -878 861 -874
rect 866 -878 878 -874
rect 885 -878 892 -874
rect 885 -881 889 -878
rect 877 -889 881 -885
rect 900 -889 904 -843
rect 912 -848 919 -844
rect 927 -850 931 -817
rect 1551 -836 1556 -807
rect 1582 -811 1586 -798
rect 1538 -841 1556 -836
rect 927 -854 995 -850
rect 927 -881 931 -854
rect 1551 -873 1556 -841
rect 1574 -815 1586 -811
rect 1604 -807 1626 -802
rect 1574 -820 1578 -815
rect 1569 -869 1574 -864
rect 1582 -873 1586 -860
rect 1604 -873 1609 -807
rect 1634 -811 1638 -798
rect 1686 -802 1690 -798
rect 1738 -802 1742 -798
rect 1626 -815 1638 -811
rect 1656 -807 1678 -802
rect 1686 -807 1730 -802
rect 1738 -807 1758 -802
rect 1626 -820 1630 -815
rect 1621 -869 1626 -864
rect 1634 -873 1638 -860
rect 1656 -873 1661 -807
rect 1675 -830 1678 -825
rect 1686 -834 1690 -807
rect 1678 -865 1682 -854
rect 1678 -869 1690 -865
rect 1551 -878 1574 -873
rect 1582 -878 1626 -873
rect 1634 -878 1678 -873
rect 1582 -881 1586 -878
rect 1634 -881 1638 -878
rect 1686 -881 1690 -869
rect 1708 -873 1713 -807
rect 1727 -830 1730 -825
rect 1738 -834 1742 -807
rect 1730 -865 1734 -854
rect 1753 -856 1758 -807
rect 1778 -804 1782 -798
rect 1810 -804 1814 -798
rect 1786 -856 1790 -844
rect 1818 -856 1822 -844
rect 1753 -861 1778 -856
rect 1786 -861 1810 -856
rect 1818 -861 1852 -856
rect 1786 -864 1790 -861
rect 1818 -864 1822 -861
rect 1730 -869 1742 -865
rect 1708 -878 1730 -873
rect 1738 -881 1742 -869
rect 907 -889 911 -885
rect 947 -889 951 -885
rect 848 -893 957 -889
rect 867 -901 909 -897
rect 1778 -891 1782 -884
rect 1810 -891 1814 -884
rect 1768 -893 1832 -891
rect 1768 -897 1770 -893
rect 1774 -897 1794 -893
rect 1798 -897 1802 -893
rect 1806 -897 1826 -893
rect 1830 -897 1832 -893
rect 1768 -899 1832 -897
rect 898 -909 929 -905
rect 1574 -909 1578 -901
rect 1626 -909 1630 -901
rect 1678 -909 1682 -901
rect 1730 -909 1734 -901
rect 1564 -910 1752 -909
rect 1564 -914 1591 -910
rect 1595 -914 1643 -910
rect 1647 -914 1695 -910
rect 1699 -914 1747 -910
rect 1751 -914 1752 -910
rect 1564 -915 1752 -914
rect 1557 -928 1564 -923
rect 1569 -928 1616 -923
rect 1621 -928 1670 -923
rect 1675 -928 1722 -923
rect 963 -974 1236 -969
rect 852 -981 880 -977
rect 852 -989 856 -981
rect 876 -989 880 -981
rect 788 -1022 856 -1018
rect 864 -1022 868 -994
rect 924 -996 948 -993
rect 930 -1002 933 -996
rect 874 -1022 925 -1021
rect 864 -1025 931 -1022
rect 939 -1022 942 -1014
rect 963 -1021 968 -974
rect 945 -1022 982 -1021
rect 939 -1025 982 -1022
rect 864 -1026 925 -1025
rect 779 -1033 868 -1029
rect 873 -1033 874 -1029
rect 779 -1034 874 -1033
rect 758 -1094 762 -1084
rect 264 -1095 762 -1094
rect 258 -1098 762 -1095
rect 183 -1099 244 -1098
rect -349 -1108 -342 -1103
rect -337 -1108 -290 -1103
rect -285 -1108 -236 -1103
rect -231 -1108 -184 -1103
rect 115 -1106 187 -1102
rect 192 -1106 193 -1102
rect 115 -1107 193 -1106
rect 196 -1110 199 -1099
rect 258 -1101 261 -1098
rect 264 -1099 762 -1098
rect 249 -1111 252 -1107
rect 243 -1114 267 -1111
rect 171 -1130 175 -1115
rect -343 -1141 -155 -1138
rect -343 -1145 -340 -1141
rect -336 -1145 -318 -1141
rect -314 -1145 -288 -1141
rect -284 -1145 -266 -1141
rect -262 -1145 -236 -1141
rect -232 -1145 -214 -1141
rect -210 -1145 -184 -1141
rect -180 -1145 -162 -1141
rect -158 -1145 -155 -1141
rect -343 -1147 -155 -1145
rect 172 -1141 200 -1137
rect -333 -1153 -329 -1147
rect -281 -1153 -277 -1147
rect -229 -1153 -225 -1147
rect -177 -1153 -173 -1147
rect 172 -1149 176 -1141
rect 196 -1149 200 -1141
rect 116 -1182 176 -1178
rect 184 -1182 188 -1154
rect 243 -1156 267 -1153
rect 249 -1162 252 -1156
rect 194 -1182 244 -1181
rect -139 -1187 -75 -1184
rect 184 -1185 250 -1182
rect 258 -1182 261 -1174
rect 315 -1177 331 -1171
rect 281 -1181 286 -1180
rect 264 -1182 291 -1181
rect 258 -1185 291 -1182
rect 184 -1186 244 -1185
rect -139 -1191 -136 -1187
rect -132 -1191 -114 -1187
rect -110 -1191 -104 -1187
rect -100 -1191 -82 -1187
rect -78 -1191 -75 -1187
rect -139 -1193 -75 -1191
rect 116 -1193 188 -1189
rect 193 -1193 194 -1189
rect -356 -1202 -333 -1197
rect -356 -1231 -351 -1202
rect -325 -1206 -321 -1193
rect -369 -1236 -351 -1231
rect -356 -1268 -351 -1236
rect -333 -1210 -321 -1206
rect -303 -1202 -281 -1197
rect -333 -1215 -329 -1210
rect -338 -1264 -333 -1259
rect -325 -1268 -321 -1255
rect -303 -1268 -298 -1202
rect -273 -1206 -269 -1193
rect -221 -1197 -217 -1193
rect -169 -1197 -165 -1193
rect -281 -1210 -269 -1206
rect -251 -1202 -229 -1197
rect -221 -1202 -177 -1197
rect -169 -1202 -149 -1197
rect -281 -1215 -277 -1210
rect -286 -1264 -281 -1259
rect -273 -1268 -269 -1255
rect -251 -1268 -246 -1202
rect -232 -1225 -229 -1220
rect -221 -1229 -217 -1202
rect -229 -1260 -225 -1249
rect -229 -1264 -217 -1260
rect -356 -1273 -333 -1268
rect -325 -1273 -281 -1268
rect -273 -1273 -229 -1268
rect -325 -1276 -321 -1273
rect -273 -1276 -269 -1273
rect -221 -1276 -217 -1264
rect -199 -1268 -194 -1202
rect -180 -1225 -177 -1220
rect -169 -1229 -165 -1202
rect -177 -1260 -173 -1249
rect -154 -1251 -149 -1202
rect -129 -1199 -125 -1193
rect -97 -1199 -93 -1193
rect 116 -1194 194 -1193
rect 197 -1197 200 -1186
rect 258 -1188 261 -1185
rect 264 -1186 291 -1185
rect 249 -1198 252 -1194
rect 243 -1201 267 -1198
rect 172 -1217 176 -1202
rect -121 -1251 -117 -1239
rect -89 -1251 -85 -1239
rect 174 -1229 202 -1225
rect 174 -1237 178 -1229
rect 198 -1237 202 -1229
rect -154 -1256 -129 -1251
rect -121 -1256 -97 -1251
rect -89 -1256 -55 -1251
rect -121 -1259 -117 -1256
rect -89 -1259 -85 -1256
rect -177 -1264 -165 -1260
rect -199 -1273 -177 -1268
rect -169 -1276 -165 -1264
rect 118 -1270 178 -1266
rect 186 -1270 190 -1242
rect 246 -1244 270 -1241
rect 252 -1250 255 -1244
rect 281 -1245 286 -1186
rect 319 -1225 328 -1177
rect 804 -1234 809 -1034
rect 816 -1125 820 -1034
rect 877 -1037 880 -1026
rect 939 -1028 942 -1025
rect 945 -1026 982 -1025
rect 930 -1038 933 -1034
rect 924 -1041 948 -1038
rect 852 -1057 856 -1042
rect 979 -1084 982 -1026
rect 1000 -1046 1034 -1043
rect 1006 -1052 1009 -1046
rect 1041 -1059 1065 -1056
rect 856 -1088 884 -1084
rect 979 -1087 1017 -1084
rect 1025 -1085 1028 -1076
rect 1047 -1065 1050 -1059
rect 856 -1096 860 -1088
rect 880 -1096 884 -1088
rect 1025 -1088 1048 -1085
rect 1056 -1085 1059 -1077
rect 1056 -1088 1076 -1085
rect 979 -1093 1007 -1090
rect 816 -1128 860 -1125
rect 816 -1129 824 -1128
rect 851 -1129 860 -1128
rect 868 -1129 872 -1101
rect 928 -1103 952 -1100
rect 934 -1109 937 -1103
rect 878 -1129 929 -1128
rect 868 -1132 935 -1129
rect 943 -1129 946 -1121
rect 979 -1126 982 -1093
rect 1025 -1091 1028 -1088
rect 1056 -1091 1059 -1088
rect 1016 -1094 1028 -1091
rect 1016 -1097 1019 -1094
rect 1047 -1101 1050 -1097
rect 1006 -1109 1009 -1103
rect 1025 -1109 1028 -1103
rect 1041 -1104 1065 -1101
rect 1000 -1112 1034 -1109
rect 949 -1129 963 -1128
rect 943 -1132 963 -1129
rect 868 -1133 929 -1132
rect 847 -1140 872 -1136
rect 877 -1140 878 -1136
rect 847 -1141 878 -1140
rect 881 -1144 884 -1133
rect 943 -1135 946 -1132
rect 949 -1133 963 -1132
rect 934 -1145 937 -1141
rect 928 -1148 952 -1145
rect 856 -1164 860 -1149
rect 1073 -1163 1076 -1088
rect 1088 -1125 1122 -1122
rect 1094 -1131 1097 -1125
rect 1129 -1138 1153 -1135
rect 1073 -1166 1105 -1163
rect 1113 -1164 1116 -1155
rect 1135 -1144 1138 -1138
rect 1113 -1167 1136 -1164
rect 1144 -1164 1147 -1156
rect 1144 -1167 1193 -1164
rect 1073 -1172 1095 -1169
rect 856 -1197 884 -1193
rect 856 -1205 860 -1197
rect 880 -1205 884 -1197
rect 804 -1238 860 -1234
rect 868 -1238 872 -1210
rect 928 -1212 952 -1209
rect 934 -1218 937 -1212
rect 1000 -1215 1034 -1212
rect 878 -1238 929 -1237
rect 868 -1241 935 -1238
rect 943 -1238 946 -1230
rect 1006 -1221 1009 -1215
rect 949 -1238 984 -1237
rect 943 -1241 985 -1238
rect 868 -1242 929 -1241
rect 281 -1249 872 -1245
rect 877 -1249 878 -1245
rect 281 -1250 878 -1249
rect 881 -1253 884 -1242
rect 943 -1244 946 -1241
rect 949 -1242 985 -1241
rect 196 -1270 247 -1269
rect 186 -1273 253 -1270
rect 261 -1270 264 -1262
rect 934 -1254 937 -1250
rect 928 -1257 952 -1254
rect 267 -1270 831 -1269
rect 261 -1273 831 -1270
rect 856 -1273 860 -1258
rect 958 -1261 963 -1242
rect 982 -1253 985 -1242
rect 1041 -1228 1065 -1225
rect 982 -1256 1017 -1253
rect 1025 -1254 1028 -1245
rect 1047 -1234 1050 -1228
rect 1025 -1257 1048 -1254
rect 1056 -1254 1059 -1246
rect 1073 -1254 1076 -1172
rect 1113 -1170 1116 -1167
rect 1144 -1170 1147 -1167
rect 1104 -1173 1116 -1170
rect 1104 -1176 1107 -1173
rect 1135 -1180 1138 -1176
rect 1094 -1188 1097 -1182
rect 1113 -1188 1116 -1182
rect 1129 -1183 1153 -1180
rect 1088 -1191 1122 -1188
rect 1056 -1257 1076 -1254
rect 973 -1262 1007 -1259
rect 186 -1274 247 -1273
rect -129 -1286 -125 -1279
rect -97 -1286 -93 -1279
rect 118 -1281 190 -1277
rect 195 -1281 196 -1277
rect 118 -1282 196 -1281
rect 199 -1285 202 -1274
rect 261 -1276 264 -1273
rect 267 -1274 831 -1273
rect -139 -1288 -75 -1286
rect -139 -1292 -137 -1288
rect -133 -1292 -113 -1288
rect -109 -1292 -105 -1288
rect -101 -1292 -81 -1288
rect -77 -1292 -75 -1288
rect -139 -1294 -75 -1292
rect 252 -1286 255 -1282
rect 246 -1289 270 -1286
rect -333 -1304 -329 -1296
rect -281 -1304 -277 -1296
rect -229 -1304 -225 -1296
rect -177 -1304 -173 -1296
rect -343 -1305 -155 -1304
rect 174 -1305 178 -1290
rect 826 -1292 831 -1274
rect 826 -1293 912 -1292
rect 973 -1293 976 -1262
rect 1025 -1260 1028 -1257
rect 1056 -1260 1059 -1257
rect 1016 -1263 1028 -1260
rect 1016 -1266 1019 -1263
rect 1047 -1270 1050 -1266
rect 1006 -1278 1009 -1272
rect 1025 -1278 1028 -1272
rect 1041 -1273 1065 -1270
rect 1000 -1281 1034 -1278
rect 826 -1296 976 -1293
rect 826 -1297 912 -1296
rect -343 -1309 -316 -1305
rect -312 -1309 -264 -1305
rect -260 -1309 -212 -1305
rect -208 -1309 -160 -1305
rect -156 -1309 -155 -1305
rect -343 -1310 -155 -1309
rect 174 -1315 202 -1311
rect -350 -1323 -343 -1318
rect -338 -1323 -291 -1318
rect -286 -1323 -237 -1318
rect -232 -1323 -185 -1318
rect 174 -1323 178 -1315
rect 198 -1323 202 -1315
rect 896 -1321 901 -1297
rect 118 -1356 178 -1352
rect 186 -1356 190 -1328
rect 247 -1330 271 -1327
rect 253 -1336 256 -1330
rect 196 -1356 248 -1355
rect 186 -1359 254 -1356
rect 262 -1356 265 -1348
rect 268 -1356 309 -1355
rect 262 -1359 309 -1356
rect 186 -1360 248 -1359
rect 118 -1367 190 -1363
rect 195 -1367 196 -1363
rect 118 -1368 196 -1367
rect -351 -1371 -163 -1368
rect 199 -1371 202 -1360
rect 262 -1362 265 -1359
rect 268 -1360 309 -1359
rect -351 -1375 -348 -1371
rect -344 -1375 -326 -1371
rect -322 -1375 -296 -1371
rect -292 -1375 -274 -1371
rect -270 -1375 -244 -1371
rect -240 -1375 -222 -1371
rect -218 -1375 -192 -1371
rect -188 -1375 -170 -1371
rect -166 -1375 -163 -1371
rect -351 -1377 -163 -1375
rect 253 -1372 256 -1368
rect 247 -1375 271 -1372
rect -341 -1383 -337 -1377
rect -289 -1383 -285 -1377
rect -237 -1383 -233 -1377
rect -185 -1383 -181 -1377
rect 174 -1391 178 -1376
rect -147 -1417 -83 -1414
rect -147 -1421 -144 -1417
rect -140 -1421 -122 -1417
rect -118 -1421 -112 -1417
rect -108 -1421 -90 -1417
rect -86 -1421 -83 -1417
rect -147 -1423 -83 -1421
rect -364 -1432 -341 -1427
rect -364 -1461 -359 -1432
rect -333 -1436 -329 -1423
rect -377 -1466 -359 -1461
rect -364 -1498 -359 -1466
rect -341 -1440 -329 -1436
rect -311 -1432 -289 -1427
rect -341 -1445 -337 -1440
rect -346 -1494 -341 -1489
rect -333 -1498 -329 -1485
rect -311 -1498 -306 -1432
rect -281 -1436 -277 -1423
rect -229 -1427 -225 -1423
rect -177 -1427 -173 -1423
rect -289 -1440 -277 -1436
rect -259 -1432 -237 -1427
rect -229 -1432 -185 -1427
rect -177 -1432 -157 -1427
rect -289 -1445 -285 -1440
rect -294 -1494 -289 -1489
rect -281 -1498 -277 -1485
rect -259 -1498 -254 -1432
rect -240 -1455 -237 -1450
rect -229 -1459 -225 -1432
rect -237 -1490 -233 -1479
rect -237 -1494 -225 -1490
rect -364 -1503 -341 -1498
rect -333 -1503 -289 -1498
rect -281 -1503 -237 -1498
rect -333 -1506 -329 -1503
rect -281 -1506 -277 -1503
rect -229 -1506 -225 -1494
rect -207 -1498 -202 -1432
rect -188 -1455 -185 -1450
rect -177 -1459 -173 -1432
rect -185 -1490 -181 -1479
rect -162 -1481 -157 -1432
rect -137 -1429 -133 -1423
rect -105 -1429 -101 -1423
rect -129 -1481 -125 -1469
rect -97 -1481 -93 -1469
rect -162 -1486 -137 -1481
rect -129 -1486 -105 -1481
rect -97 -1486 -63 -1481
rect -129 -1489 -125 -1486
rect -97 -1489 -93 -1486
rect -185 -1494 -173 -1490
rect -207 -1503 -185 -1498
rect -177 -1506 -173 -1494
rect -137 -1516 -133 -1509
rect -105 -1516 -101 -1509
rect -147 -1518 -83 -1516
rect -147 -1522 -145 -1518
rect -141 -1522 -121 -1518
rect -117 -1522 -113 -1518
rect -109 -1522 -89 -1518
rect -85 -1522 -83 -1518
rect -147 -1524 -83 -1522
rect -341 -1534 -337 -1526
rect -289 -1534 -285 -1526
rect -237 -1534 -233 -1526
rect -185 -1534 -181 -1526
rect -351 -1535 -163 -1534
rect -351 -1539 -324 -1535
rect -320 -1539 -272 -1535
rect -268 -1539 -220 -1535
rect -216 -1539 -168 -1535
rect -164 -1539 -163 -1535
rect -351 -1540 -163 -1539
rect -358 -1553 -351 -1548
rect -346 -1553 -299 -1548
rect -294 -1553 -245 -1548
rect -240 -1553 -193 -1548
rect -349 -1597 -161 -1594
rect -349 -1601 -346 -1597
rect -342 -1601 -324 -1597
rect -320 -1601 -294 -1597
rect -290 -1601 -272 -1597
rect -268 -1601 -242 -1597
rect -238 -1601 -220 -1597
rect -216 -1601 -190 -1597
rect -186 -1601 -168 -1597
rect -164 -1601 -161 -1597
rect -349 -1603 -161 -1601
rect -339 -1609 -335 -1603
rect -287 -1609 -283 -1603
rect -235 -1609 -231 -1603
rect -183 -1609 -179 -1603
rect -145 -1643 -81 -1640
rect -145 -1647 -142 -1643
rect -138 -1647 -120 -1643
rect -116 -1647 -110 -1643
rect -106 -1647 -88 -1643
rect -84 -1647 -81 -1643
rect -145 -1649 -81 -1647
rect -362 -1658 -339 -1653
rect -362 -1687 -357 -1658
rect -331 -1662 -327 -1649
rect -375 -1692 -357 -1687
rect -362 -1724 -357 -1692
rect -339 -1666 -327 -1662
rect -309 -1658 -287 -1653
rect -339 -1671 -335 -1666
rect -344 -1720 -339 -1715
rect -331 -1724 -327 -1711
rect -309 -1724 -304 -1658
rect -279 -1662 -275 -1649
rect -227 -1653 -223 -1649
rect -175 -1653 -171 -1649
rect -287 -1666 -275 -1662
rect -257 -1658 -235 -1653
rect -227 -1658 -183 -1653
rect -175 -1658 -155 -1653
rect -287 -1671 -283 -1666
rect -292 -1720 -287 -1715
rect -279 -1724 -275 -1711
rect -257 -1724 -252 -1658
rect -238 -1681 -235 -1676
rect -227 -1685 -223 -1658
rect -235 -1716 -231 -1705
rect -235 -1720 -223 -1716
rect -362 -1729 -339 -1724
rect -331 -1729 -287 -1724
rect -279 -1729 -235 -1724
rect -331 -1732 -327 -1729
rect -279 -1732 -275 -1729
rect -227 -1732 -223 -1720
rect -205 -1724 -200 -1658
rect -186 -1681 -183 -1676
rect -175 -1685 -171 -1658
rect -183 -1716 -179 -1705
rect -160 -1707 -155 -1658
rect -135 -1655 -131 -1649
rect -103 -1655 -99 -1649
rect -127 -1707 -123 -1695
rect -95 -1707 -91 -1695
rect -160 -1712 -135 -1707
rect -127 -1712 -103 -1707
rect -95 -1712 -61 -1707
rect -127 -1715 -123 -1712
rect -95 -1715 -91 -1712
rect -183 -1720 -171 -1716
rect -205 -1729 -183 -1724
rect -175 -1732 -171 -1720
rect -135 -1742 -131 -1735
rect -103 -1742 -99 -1735
rect -145 -1744 -81 -1742
rect -145 -1748 -143 -1744
rect -139 -1748 -119 -1744
rect -115 -1748 -111 -1744
rect -107 -1748 -87 -1744
rect -83 -1748 -81 -1744
rect -145 -1750 -81 -1748
rect -339 -1760 -335 -1752
rect -287 -1760 -283 -1752
rect -235 -1760 -231 -1752
rect -183 -1760 -179 -1752
rect -349 -1761 -161 -1760
rect -349 -1765 -322 -1761
rect -318 -1765 -270 -1761
rect -266 -1765 -218 -1761
rect -214 -1765 -166 -1761
rect -162 -1765 -161 -1761
rect -349 -1766 -161 -1765
rect -356 -1779 -349 -1774
rect -344 -1779 -297 -1774
rect -292 -1779 -243 -1774
rect -238 -1779 -191 -1774
rect -349 -1820 -161 -1817
rect -349 -1824 -346 -1820
rect -342 -1824 -324 -1820
rect -320 -1824 -294 -1820
rect -290 -1824 -272 -1820
rect -268 -1824 -242 -1820
rect -238 -1824 -220 -1820
rect -216 -1824 -190 -1820
rect -186 -1824 -168 -1820
rect -164 -1824 -161 -1820
rect -349 -1826 -161 -1824
rect -339 -1832 -335 -1826
rect -287 -1832 -283 -1826
rect -235 -1832 -231 -1826
rect -183 -1832 -179 -1826
rect 302 -1827 307 -1360
rect 349 -1354 378 -1353
rect 343 -1355 380 -1354
rect 343 -1360 1169 -1355
rect 936 -1668 941 -1360
rect 1164 -1460 1169 -1360
rect 1231 -1449 1236 -974
rect 1564 -979 1752 -976
rect 1564 -983 1567 -979
rect 1571 -983 1589 -979
rect 1593 -983 1619 -979
rect 1623 -983 1641 -979
rect 1645 -983 1671 -979
rect 1675 -983 1693 -979
rect 1697 -983 1723 -979
rect 1727 -983 1745 -979
rect 1749 -983 1752 -979
rect 1564 -985 1752 -983
rect 1574 -991 1578 -985
rect 1626 -991 1630 -985
rect 1678 -991 1682 -985
rect 1730 -991 1734 -985
rect 1768 -1025 1832 -1022
rect 1768 -1029 1771 -1025
rect 1775 -1029 1793 -1025
rect 1797 -1029 1803 -1025
rect 1807 -1029 1825 -1025
rect 1829 -1029 1832 -1025
rect 1768 -1031 1832 -1029
rect 1551 -1040 1574 -1035
rect 1551 -1069 1556 -1040
rect 1582 -1044 1586 -1031
rect 1538 -1074 1556 -1069
rect 1292 -1089 1401 -1085
rect 1273 -1104 1283 -1100
rect 1279 -1110 1283 -1104
rect 1279 -1114 1296 -1110
rect 1306 -1135 1310 -1089
rect 1321 -1095 1325 -1089
rect 1351 -1095 1355 -1089
rect 1391 -1095 1395 -1089
rect 1329 -1110 1333 -1103
rect 1318 -1114 1322 -1110
rect 1329 -1114 1353 -1110
rect 1329 -1117 1333 -1114
rect 1321 -1125 1325 -1121
rect 1315 -1129 1348 -1125
rect 1306 -1139 1339 -1135
rect 1321 -1145 1325 -1139
rect 1329 -1160 1333 -1153
rect 1286 -1164 1305 -1160
rect 1310 -1164 1322 -1160
rect 1329 -1164 1336 -1160
rect 1329 -1167 1333 -1164
rect 1321 -1175 1325 -1171
rect 1344 -1175 1348 -1129
rect 1356 -1134 1363 -1130
rect 1371 -1136 1375 -1103
rect 1551 -1106 1556 -1074
rect 1574 -1048 1586 -1044
rect 1604 -1040 1626 -1035
rect 1574 -1053 1578 -1048
rect 1569 -1102 1574 -1097
rect 1582 -1106 1586 -1093
rect 1604 -1106 1609 -1040
rect 1634 -1044 1638 -1031
rect 1686 -1035 1690 -1031
rect 1738 -1035 1742 -1031
rect 1626 -1048 1638 -1044
rect 1656 -1040 1678 -1035
rect 1686 -1040 1730 -1035
rect 1738 -1040 1758 -1035
rect 1626 -1053 1630 -1048
rect 1621 -1102 1626 -1097
rect 1634 -1106 1638 -1093
rect 1656 -1106 1661 -1040
rect 1675 -1063 1678 -1058
rect 1686 -1067 1690 -1040
rect 1678 -1098 1682 -1087
rect 1678 -1102 1690 -1098
rect 1551 -1111 1574 -1106
rect 1582 -1111 1626 -1106
rect 1634 -1111 1678 -1106
rect 1582 -1114 1586 -1111
rect 1634 -1114 1638 -1111
rect 1686 -1114 1690 -1102
rect 1708 -1106 1713 -1040
rect 1727 -1063 1730 -1058
rect 1738 -1067 1742 -1040
rect 1730 -1098 1734 -1087
rect 1753 -1089 1758 -1040
rect 1778 -1037 1782 -1031
rect 1810 -1037 1814 -1031
rect 1786 -1089 1790 -1077
rect 1818 -1089 1822 -1077
rect 1753 -1094 1778 -1089
rect 1786 -1094 1810 -1089
rect 1818 -1094 1852 -1089
rect 1786 -1097 1790 -1094
rect 1818 -1097 1822 -1094
rect 1730 -1102 1742 -1098
rect 1708 -1111 1730 -1106
rect 1738 -1114 1742 -1102
rect 1778 -1124 1782 -1117
rect 1810 -1124 1814 -1117
rect 1768 -1126 1832 -1124
rect 1768 -1130 1770 -1126
rect 1774 -1130 1794 -1126
rect 1798 -1130 1802 -1126
rect 1806 -1130 1826 -1126
rect 1830 -1130 1832 -1126
rect 1768 -1132 1832 -1130
rect 1371 -1140 1452 -1136
rect 1371 -1167 1375 -1140
rect 1574 -1142 1578 -1134
rect 1626 -1142 1630 -1134
rect 1678 -1142 1682 -1134
rect 1730 -1142 1734 -1134
rect 1564 -1143 1752 -1142
rect 1564 -1147 1591 -1143
rect 1595 -1147 1643 -1143
rect 1647 -1147 1695 -1143
rect 1699 -1147 1747 -1143
rect 1751 -1147 1752 -1143
rect 1564 -1148 1752 -1147
rect 1557 -1161 1564 -1156
rect 1569 -1161 1616 -1156
rect 1621 -1161 1670 -1156
rect 1675 -1161 1722 -1156
rect 1351 -1175 1355 -1171
rect 1391 -1175 1395 -1171
rect 1292 -1179 1401 -1175
rect 1311 -1187 1353 -1183
rect 1342 -1195 1373 -1191
rect 1559 -1205 1747 -1202
rect 1559 -1209 1562 -1205
rect 1566 -1209 1584 -1205
rect 1588 -1209 1614 -1205
rect 1618 -1209 1636 -1205
rect 1640 -1209 1666 -1205
rect 1670 -1209 1688 -1205
rect 1692 -1209 1718 -1205
rect 1722 -1209 1740 -1205
rect 1744 -1209 1747 -1205
rect 1559 -1211 1747 -1209
rect 1569 -1217 1573 -1211
rect 1621 -1217 1625 -1211
rect 1673 -1217 1677 -1211
rect 1725 -1217 1729 -1211
rect 1763 -1251 1827 -1248
rect 1763 -1255 1766 -1251
rect 1770 -1255 1788 -1251
rect 1792 -1255 1798 -1251
rect 1802 -1255 1820 -1251
rect 1824 -1255 1827 -1251
rect 1763 -1257 1827 -1255
rect 1546 -1266 1569 -1261
rect 1546 -1295 1551 -1266
rect 1577 -1270 1581 -1257
rect 1533 -1300 1551 -1295
rect 1546 -1332 1551 -1300
rect 1569 -1274 1581 -1270
rect 1599 -1266 1621 -1261
rect 1569 -1279 1573 -1274
rect 1564 -1328 1569 -1323
rect 1577 -1332 1581 -1319
rect 1599 -1332 1604 -1266
rect 1629 -1270 1633 -1257
rect 1681 -1261 1685 -1257
rect 1733 -1261 1737 -1257
rect 1621 -1274 1633 -1270
rect 1651 -1266 1673 -1261
rect 1681 -1266 1725 -1261
rect 1733 -1266 1753 -1261
rect 1621 -1279 1625 -1274
rect 1616 -1328 1621 -1323
rect 1629 -1332 1633 -1319
rect 1651 -1332 1656 -1266
rect 1670 -1289 1673 -1284
rect 1681 -1293 1685 -1266
rect 1673 -1324 1677 -1313
rect 1673 -1328 1685 -1324
rect 1546 -1337 1569 -1332
rect 1577 -1337 1621 -1332
rect 1629 -1337 1673 -1332
rect 1577 -1340 1581 -1337
rect 1629 -1340 1633 -1337
rect 1681 -1340 1685 -1328
rect 1703 -1332 1708 -1266
rect 1722 -1289 1725 -1284
rect 1733 -1293 1737 -1266
rect 1725 -1324 1729 -1313
rect 1748 -1315 1753 -1266
rect 1773 -1263 1777 -1257
rect 1805 -1263 1809 -1257
rect 1781 -1315 1785 -1303
rect 1813 -1315 1817 -1303
rect 1748 -1320 1773 -1315
rect 1781 -1320 1805 -1315
rect 1813 -1320 1847 -1315
rect 1781 -1323 1785 -1320
rect 1813 -1323 1817 -1320
rect 1725 -1328 1737 -1324
rect 1703 -1337 1725 -1332
rect 1733 -1340 1737 -1328
rect 1773 -1350 1777 -1343
rect 1805 -1350 1809 -1343
rect 1763 -1352 1827 -1350
rect 1763 -1356 1765 -1352
rect 1769 -1356 1789 -1352
rect 1793 -1356 1797 -1352
rect 1801 -1356 1821 -1352
rect 1825 -1356 1827 -1352
rect 1763 -1358 1827 -1356
rect 1569 -1368 1573 -1360
rect 1621 -1368 1625 -1360
rect 1673 -1368 1677 -1360
rect 1725 -1368 1729 -1360
rect 1559 -1369 1747 -1368
rect 1559 -1373 1586 -1369
rect 1590 -1373 1638 -1369
rect 1642 -1373 1690 -1369
rect 1694 -1373 1742 -1369
rect 1746 -1373 1747 -1369
rect 1559 -1374 1747 -1373
rect 1552 -1387 1559 -1382
rect 1564 -1387 1611 -1382
rect 1616 -1387 1665 -1382
rect 1670 -1387 1717 -1382
rect 1256 -1412 1284 -1408
rect 1256 -1420 1260 -1412
rect 1280 -1420 1284 -1412
rect 1231 -1453 1260 -1449
rect 1268 -1453 1272 -1425
rect 1328 -1427 1352 -1424
rect 1334 -1433 1337 -1427
rect 1278 -1453 1329 -1452
rect 1268 -1456 1335 -1453
rect 1343 -1453 1346 -1445
rect 1349 -1453 1360 -1452
rect 1343 -1456 1367 -1453
rect 1268 -1457 1329 -1456
rect 1164 -1464 1272 -1460
rect 1277 -1464 1278 -1460
rect 1164 -1465 1278 -1464
rect 1195 -1565 1200 -1465
rect 1281 -1468 1284 -1457
rect 1343 -1459 1346 -1456
rect 1349 -1457 1360 -1456
rect 1334 -1469 1337 -1465
rect 1328 -1472 1352 -1469
rect 1256 -1488 1260 -1473
rect 1364 -1502 1367 -1456
rect 1388 -1464 1422 -1461
rect 1394 -1470 1397 -1464
rect 1429 -1477 1453 -1474
rect 1364 -1505 1405 -1502
rect 1413 -1503 1416 -1494
rect 1435 -1483 1438 -1477
rect 1413 -1506 1436 -1503
rect 1444 -1503 1447 -1495
rect 1444 -1506 1493 -1503
rect 1371 -1511 1395 -1508
rect 1256 -1517 1284 -1513
rect 1256 -1525 1260 -1517
rect 1280 -1525 1284 -1517
rect 1241 -1558 1260 -1554
rect 1268 -1558 1272 -1530
rect 1328 -1532 1352 -1529
rect 1334 -1538 1337 -1532
rect 1278 -1558 1329 -1557
rect 1268 -1561 1335 -1558
rect 1343 -1558 1346 -1550
rect 1349 -1558 1360 -1557
rect 1371 -1558 1374 -1511
rect 1413 -1509 1416 -1506
rect 1444 -1509 1447 -1506
rect 1404 -1512 1416 -1509
rect 1404 -1515 1407 -1512
rect 1435 -1519 1438 -1515
rect 1394 -1527 1397 -1521
rect 1413 -1527 1416 -1521
rect 1429 -1522 1453 -1519
rect 1388 -1530 1422 -1527
rect 1343 -1561 1374 -1558
rect 1268 -1562 1329 -1561
rect 1195 -1569 1272 -1565
rect 1277 -1569 1278 -1565
rect 1195 -1570 1278 -1569
rect 1281 -1573 1284 -1562
rect 1343 -1564 1346 -1561
rect 1349 -1562 1360 -1561
rect 1334 -1574 1337 -1570
rect 1328 -1577 1352 -1574
rect 1256 -1593 1260 -1578
rect 1487 -1615 1490 -1506
rect 1501 -1577 1535 -1574
rect 1507 -1583 1510 -1577
rect 1542 -1590 1566 -1587
rect 1256 -1620 1284 -1616
rect 1487 -1618 1518 -1615
rect 1526 -1616 1529 -1607
rect 1548 -1596 1551 -1590
rect 1256 -1628 1260 -1620
rect 1280 -1628 1284 -1620
rect 1526 -1619 1549 -1616
rect 1557 -1616 1560 -1608
rect 1557 -1619 1597 -1616
rect 1488 -1624 1508 -1621
rect 1250 -1661 1260 -1657
rect 1268 -1661 1272 -1633
rect 1328 -1635 1352 -1632
rect 1334 -1641 1337 -1635
rect 1278 -1661 1329 -1660
rect 1268 -1664 1335 -1661
rect 1343 -1661 1346 -1653
rect 1349 -1661 1360 -1660
rect 1343 -1664 1369 -1661
rect 1268 -1665 1329 -1664
rect 936 -1672 1272 -1668
rect 1277 -1672 1278 -1668
rect 936 -1673 1278 -1672
rect 1123 -1746 1127 -1673
rect 1281 -1676 1284 -1665
rect 1343 -1667 1346 -1664
rect 1349 -1665 1360 -1664
rect 1334 -1677 1337 -1673
rect 1328 -1680 1352 -1677
rect 1256 -1696 1260 -1681
rect 1366 -1704 1369 -1664
rect 1385 -1666 1419 -1663
rect 1391 -1672 1394 -1666
rect 1426 -1679 1450 -1676
rect 1246 -1709 1274 -1705
rect 1366 -1707 1402 -1704
rect 1410 -1705 1413 -1696
rect 1432 -1685 1435 -1679
rect 1246 -1717 1250 -1709
rect 1270 -1717 1274 -1709
rect 1410 -1708 1433 -1705
rect 1441 -1705 1444 -1697
rect 1488 -1705 1491 -1624
rect 1526 -1622 1529 -1619
rect 1557 -1622 1560 -1619
rect 1517 -1625 1529 -1622
rect 1517 -1628 1520 -1625
rect 1548 -1632 1551 -1628
rect 1507 -1640 1510 -1634
rect 1526 -1640 1529 -1634
rect 1542 -1635 1566 -1632
rect 1501 -1643 1535 -1640
rect 1441 -1708 1494 -1705
rect 1358 -1713 1392 -1710
rect 1123 -1750 1250 -1746
rect 1258 -1750 1262 -1722
rect 1318 -1724 1342 -1721
rect 1324 -1730 1327 -1724
rect 1268 -1750 1319 -1749
rect 1258 -1753 1325 -1750
rect 1333 -1750 1336 -1742
rect 1358 -1749 1361 -1713
rect 1410 -1711 1413 -1708
rect 1441 -1711 1444 -1708
rect 1401 -1714 1413 -1711
rect 1401 -1717 1404 -1714
rect 1594 -1717 1597 -1619
rect 1604 -1679 1638 -1676
rect 1610 -1685 1613 -1679
rect 1645 -1692 1669 -1689
rect 1432 -1721 1435 -1717
rect 1594 -1720 1621 -1717
rect 1629 -1718 1632 -1709
rect 1651 -1698 1654 -1692
rect 1629 -1721 1652 -1718
rect 1660 -1718 1663 -1710
rect 1660 -1721 1723 -1718
rect 1391 -1729 1394 -1723
rect 1410 -1729 1413 -1723
rect 1426 -1724 1450 -1721
rect 1587 -1726 1611 -1723
rect 1385 -1732 1419 -1729
rect 1339 -1750 1361 -1749
rect 1333 -1752 1361 -1750
rect 1333 -1753 1350 -1752
rect 1258 -1754 1319 -1753
rect 1238 -1761 1262 -1757
rect 1267 -1761 1268 -1757
rect 1238 -1762 1268 -1761
rect 1238 -1764 1241 -1762
rect 1271 -1765 1274 -1754
rect 1333 -1756 1336 -1753
rect 1339 -1754 1350 -1753
rect 1324 -1766 1327 -1762
rect 1318 -1769 1342 -1766
rect 1246 -1785 1250 -1770
rect 1587 -1827 1590 -1726
rect 1629 -1724 1632 -1721
rect 1660 -1724 1663 -1721
rect 1620 -1727 1632 -1724
rect 1620 -1730 1623 -1727
rect 1651 -1734 1654 -1730
rect 1610 -1742 1613 -1736
rect 1629 -1742 1632 -1736
rect 1645 -1737 1669 -1734
rect 1604 -1745 1638 -1742
rect 302 -1832 1595 -1827
rect -145 -1866 -81 -1863
rect -145 -1870 -142 -1866
rect -138 -1870 -120 -1866
rect -116 -1870 -110 -1866
rect -106 -1870 -88 -1866
rect -84 -1870 -81 -1866
rect -145 -1872 -81 -1870
rect -362 -1881 -339 -1876
rect -362 -1910 -357 -1881
rect -331 -1885 -327 -1872
rect -375 -1915 -357 -1910
rect -362 -1947 -357 -1915
rect -339 -1889 -327 -1885
rect -309 -1881 -287 -1876
rect -339 -1894 -335 -1889
rect -344 -1943 -339 -1938
rect -331 -1947 -327 -1934
rect -309 -1947 -304 -1881
rect -279 -1885 -275 -1872
rect -227 -1876 -223 -1872
rect -175 -1876 -171 -1872
rect -287 -1889 -275 -1885
rect -257 -1881 -235 -1876
rect -227 -1881 -183 -1876
rect -175 -1881 -155 -1876
rect -287 -1894 -283 -1889
rect -292 -1943 -287 -1938
rect -279 -1947 -275 -1934
rect -257 -1947 -252 -1881
rect -238 -1904 -235 -1899
rect -227 -1908 -223 -1881
rect -235 -1939 -231 -1928
rect -235 -1943 -223 -1939
rect -362 -1952 -339 -1947
rect -331 -1952 -287 -1947
rect -279 -1952 -235 -1947
rect -331 -1955 -327 -1952
rect -279 -1955 -275 -1952
rect -227 -1955 -223 -1943
rect -205 -1947 -200 -1881
rect -186 -1904 -183 -1899
rect -175 -1908 -171 -1881
rect -183 -1939 -179 -1928
rect -160 -1930 -155 -1881
rect -135 -1878 -131 -1872
rect -103 -1878 -99 -1872
rect -127 -1930 -123 -1918
rect -95 -1930 -91 -1918
rect -160 -1935 -135 -1930
rect -127 -1935 -103 -1930
rect -95 -1935 -61 -1930
rect -127 -1938 -123 -1935
rect -95 -1938 -91 -1935
rect -183 -1943 -171 -1939
rect -205 -1952 -183 -1947
rect -175 -1955 -171 -1943
rect -135 -1965 -131 -1958
rect -103 -1965 -99 -1958
rect -145 -1967 -81 -1965
rect -145 -1971 -143 -1967
rect -139 -1971 -119 -1967
rect -115 -1971 -111 -1967
rect -107 -1971 -87 -1967
rect -83 -1971 -81 -1967
rect -145 -1973 -81 -1971
rect -339 -1983 -335 -1975
rect -287 -1983 -283 -1975
rect -235 -1983 -231 -1975
rect -183 -1983 -179 -1975
rect -349 -1984 -161 -1983
rect -349 -1988 -322 -1984
rect -318 -1988 -270 -1984
rect -266 -1988 -218 -1984
rect -214 -1988 -166 -1984
rect -162 -1988 -161 -1984
rect -349 -1989 -161 -1988
rect -356 -2002 -349 -1997
rect -344 -2002 -297 -1997
rect -292 -2002 -243 -1997
rect -238 -2002 -191 -1997
<< m2contact >>
rect -336 -377 -331 -372
rect -284 -377 -279 -372
rect -230 -338 -225 -333
rect -178 -338 -173 -333
rect 1571 -391 1576 -386
rect 1623 -391 1628 -386
rect 1677 -352 1682 -347
rect 1729 -352 1734 -347
rect -336 -436 -331 -431
rect -284 -436 -279 -431
rect -230 -436 -225 -431
rect -178 -436 -173 -431
rect 1571 -450 1576 -445
rect 1623 -450 1628 -445
rect 1677 -450 1682 -445
rect 1729 -450 1734 -445
rect 125 -481 130 -476
rect 142 -481 147 -476
rect 134 -531 139 -526
rect 165 -531 170 -526
rect -339 -604 -334 -599
rect -287 -604 -282 -599
rect -233 -565 -228 -560
rect -181 -565 -176 -560
rect 180 -501 185 -496
rect 135 -553 140 -548
rect 166 -561 171 -556
rect 126 -602 131 -597
rect 143 -602 148 -597
rect 135 -652 140 -647
rect 166 -652 171 -647
rect -339 -663 -334 -658
rect -287 -663 -282 -658
rect -233 -663 -228 -658
rect -181 -663 -176 -658
rect 181 -622 186 -617
rect 368 -616 386 -598
rect 136 -674 141 -669
rect 167 -682 172 -677
rect 317 -693 334 -677
rect 126 -723 131 -718
rect 143 -723 148 -718
rect -342 -833 -337 -828
rect -290 -833 -285 -828
rect -236 -794 -231 -789
rect -184 -794 -179 -789
rect 135 -773 140 -768
rect 166 -773 171 -768
rect 181 -743 186 -738
rect 136 -795 141 -790
rect 167 -803 172 -798
rect 126 -843 131 -838
rect 143 -843 148 -838
rect -342 -892 -337 -887
rect -290 -892 -285 -887
rect -236 -892 -231 -887
rect -184 -892 -179 -887
rect 135 -893 140 -888
rect 166 -893 171 -888
rect 181 -863 186 -858
rect 136 -915 141 -910
rect 167 -923 172 -918
rect -342 -1049 -337 -1044
rect -290 -1049 -285 -1044
rect -236 -1010 -231 -1005
rect -184 -1010 -179 -1005
rect 332 -1004 352 -985
rect 563 -564 583 -550
rect 862 -570 885 -550
rect 938 -551 943 -546
rect 955 -551 960 -546
rect 947 -601 952 -596
rect 978 -601 983 -596
rect 993 -571 998 -566
rect 948 -623 953 -618
rect 979 -631 984 -626
rect 1563 -633 1568 -628
rect 1615 -633 1620 -628
rect 1669 -594 1674 -589
rect 1721 -594 1726 -589
rect 730 -729 750 -717
rect 361 -1039 378 -1021
rect 317 -1087 338 -1071
rect 528 -1059 545 -1047
rect 723 -895 736 -885
rect 549 -1089 566 -1074
rect 780 -734 798 -714
rect 918 -680 938 -662
rect 948 -675 953 -670
rect 965 -675 970 -670
rect 957 -725 962 -720
rect 988 -725 993 -720
rect 1003 -695 1008 -690
rect 1563 -692 1568 -687
rect 1615 -692 1620 -687
rect 1669 -692 1674 -687
rect 1721 -692 1726 -687
rect 958 -747 963 -742
rect 989 -755 994 -750
rect 806 -850 839 -814
rect 852 -829 857 -824
rect 869 -829 874 -824
rect 817 -879 838 -869
rect 861 -879 866 -874
rect 892 -879 897 -874
rect 907 -849 912 -844
rect 1564 -869 1569 -864
rect 1616 -869 1621 -864
rect 1670 -830 1675 -825
rect 1722 -830 1727 -825
rect 862 -901 867 -896
rect 893 -909 898 -904
rect 1564 -928 1569 -923
rect 1616 -928 1621 -923
rect 1670 -928 1675 -923
rect 1722 -928 1727 -923
rect 767 -1036 779 -1022
rect -342 -1108 -337 -1103
rect -290 -1108 -285 -1103
rect -236 -1108 -231 -1103
rect -184 -1108 -179 -1103
rect 311 -1171 336 -1150
rect -343 -1264 -338 -1259
rect -291 -1264 -286 -1259
rect -237 -1225 -232 -1220
rect -185 -1225 -180 -1220
rect 291 -1194 306 -1177
rect 318 -1238 334 -1225
rect 829 -1145 847 -1131
rect 963 -1139 983 -1126
rect 1193 -1173 1211 -1156
rect 952 -1273 967 -1261
rect -343 -1323 -338 -1318
rect -291 -1323 -286 -1318
rect -237 -1323 -232 -1318
rect -185 -1323 -180 -1318
rect -351 -1494 -346 -1489
rect -299 -1494 -294 -1489
rect -245 -1455 -240 -1450
rect -193 -1455 -188 -1450
rect -351 -1553 -346 -1548
rect -299 -1553 -294 -1548
rect -245 -1553 -240 -1548
rect -193 -1553 -188 -1548
rect -349 -1720 -344 -1715
rect -297 -1720 -292 -1715
rect -243 -1681 -238 -1676
rect -191 -1681 -186 -1676
rect -349 -1779 -344 -1774
rect -297 -1779 -292 -1774
rect -243 -1779 -238 -1774
rect -191 -1779 -186 -1774
rect 319 -1369 343 -1342
rect 889 -1345 920 -1321
rect 1251 -1112 1273 -1088
rect 1296 -1115 1301 -1110
rect 1313 -1115 1318 -1110
rect 1264 -1171 1286 -1156
rect 1305 -1165 1310 -1160
rect 1336 -1165 1341 -1160
rect 1351 -1135 1356 -1130
rect 1564 -1102 1569 -1097
rect 1616 -1102 1621 -1097
rect 1670 -1063 1675 -1058
rect 1722 -1063 1727 -1058
rect 1564 -1161 1569 -1156
rect 1616 -1161 1621 -1156
rect 1670 -1161 1675 -1156
rect 1722 -1161 1727 -1156
rect 1306 -1187 1311 -1182
rect 1337 -1195 1342 -1190
rect 1559 -1328 1564 -1323
rect 1611 -1328 1616 -1323
rect 1665 -1289 1670 -1284
rect 1717 -1289 1722 -1284
rect 1559 -1387 1564 -1382
rect 1611 -1387 1616 -1382
rect 1665 -1387 1670 -1382
rect 1717 -1387 1722 -1382
rect 1210 -1560 1241 -1536
rect 1225 -1665 1250 -1645
rect 1224 -1765 1238 -1753
rect -349 -1943 -344 -1938
rect -297 -1943 -292 -1938
rect -243 -1904 -238 -1899
rect -191 -1904 -186 -1899
rect -349 -2002 -344 -1997
rect -297 -2002 -292 -1997
rect -243 -2002 -238 -1997
rect -191 -2002 -186 -1997
<< metal2 >>
rect -336 -431 -331 -377
rect -284 -431 -279 -377
rect -230 -431 -225 -338
rect -178 -431 -173 -338
rect 1571 -445 1576 -391
rect 1623 -445 1628 -391
rect 1677 -445 1682 -352
rect 1729 -445 1734 -352
rect 130 -481 142 -477
rect 126 -496 130 -481
rect 126 -500 180 -496
rect 135 -548 139 -531
rect 166 -556 170 -531
rect -339 -658 -334 -604
rect -287 -658 -282 -604
rect -233 -658 -228 -565
rect 583 -562 862 -555
rect -181 -658 -176 -565
rect 943 -551 955 -547
rect 939 -566 943 -551
rect 939 -570 993 -566
rect 131 -602 143 -598
rect 127 -617 131 -602
rect 386 -604 871 -598
rect 127 -621 181 -617
rect 865 -634 871 -604
rect 948 -618 952 -601
rect 979 -626 983 -601
rect 865 -640 926 -634
rect 136 -669 140 -652
rect 167 -677 171 -652
rect 920 -662 926 -640
rect 953 -675 965 -671
rect 334 -691 596 -683
rect 588 -706 596 -691
rect 949 -690 953 -675
rect 1563 -687 1568 -633
rect 949 -694 1003 -690
rect 1615 -687 1620 -633
rect 1669 -687 1674 -594
rect 1721 -687 1726 -594
rect 684 -705 819 -697
rect 684 -706 692 -705
rect 588 -714 692 -706
rect 131 -723 143 -719
rect 127 -738 131 -723
rect 750 -726 780 -719
rect 127 -742 181 -738
rect -342 -887 -337 -833
rect -290 -887 -285 -833
rect -236 -887 -231 -794
rect -184 -887 -179 -794
rect 136 -790 140 -773
rect 167 -798 171 -773
rect 811 -814 819 -705
rect 958 -742 962 -725
rect 989 -750 993 -725
rect 131 -843 143 -839
rect 127 -858 131 -843
rect 857 -829 869 -825
rect 853 -844 857 -829
rect 853 -848 907 -844
rect 127 -862 181 -858
rect 136 -910 140 -893
rect 167 -918 171 -893
rect 818 -888 822 -879
rect 736 -892 822 -888
rect 862 -896 866 -879
rect 893 -904 897 -879
rect 1564 -923 1569 -869
rect 1616 -923 1621 -869
rect 1670 -923 1675 -830
rect 1722 -923 1727 -830
rect 801 -939 1260 -934
rect 352 -991 357 -988
rect 801 -991 806 -939
rect 352 -996 806 -991
rect 352 -998 357 -996
rect -342 -1103 -337 -1049
rect -290 -1103 -285 -1049
rect -236 -1103 -231 -1010
rect -184 -1103 -179 -1010
rect 378 -1033 767 -1025
rect 545 -1056 789 -1049
rect 319 -1150 328 -1087
rect 553 -1181 558 -1089
rect 782 -1134 789 -1056
rect 1255 -1088 1260 -939
rect 1301 -1115 1313 -1111
rect 782 -1141 829 -1134
rect 1297 -1130 1301 -1115
rect 1297 -1134 1351 -1130
rect 969 -1143 979 -1139
rect 306 -1186 558 -1181
rect 970 -1199 974 -1143
rect 1564 -1156 1569 -1102
rect 1211 -1167 1264 -1162
rect 1616 -1156 1621 -1102
rect 1670 -1156 1675 -1063
rect 1722 -1156 1727 -1063
rect 1306 -1182 1310 -1165
rect 1337 -1190 1341 -1165
rect 970 -1203 1218 -1199
rect -343 -1318 -338 -1264
rect -291 -1318 -286 -1264
rect -237 -1318 -232 -1225
rect -185 -1318 -180 -1225
rect 320 -1342 330 -1238
rect -351 -1548 -346 -1494
rect -299 -1548 -294 -1494
rect -245 -1548 -240 -1455
rect -193 -1548 -188 -1455
rect -349 -1774 -344 -1720
rect -297 -1774 -292 -1720
rect -243 -1774 -238 -1681
rect -191 -1774 -186 -1681
rect 892 -1753 904 -1345
rect 955 -1392 964 -1273
rect 955 -1401 1155 -1392
rect 1146 -1655 1155 -1401
rect 1214 -1536 1218 -1203
rect 1559 -1382 1564 -1328
rect 1611 -1382 1616 -1328
rect 1665 -1382 1670 -1289
rect 1717 -1382 1722 -1289
rect 1146 -1664 1225 -1655
rect 892 -1765 1224 -1753
rect -349 -1997 -344 -1943
rect -297 -1997 -292 -1943
rect -243 -1997 -238 -1904
rect -191 -1997 -186 -1904
<< labels >>
rlabel metal1 121 -455 230 -451 5 vdd
rlabel metal1 121 -545 230 -541 1 gnd
rlabel metal1 16 -478 40 -478 1 a0
rlabel metal1 15 -528 39 -528 1 b0
rlabel metal1 253 -504 278 -504 1 p0
rlabel metal1 122 -576 231 -572 5 vdd
rlabel metal1 122 -666 231 -662 1 gnd
rlabel metal1 19 -599 39 -599 1 a1
rlabel metal1 27 -649 27 -649 1 b1
rlabel metal1 267 -625 267 -625 1 p1
rlabel metal1 122 -697 231 -693 5 vdd
rlabel metal1 122 -787 231 -783 1 gnd
rlabel metal1 29 -720 29 -720 1 a2
rlabel metal1 27 -771 27 -770 1 b2
rlabel metal1 267 -746 267 -746 1 p2
rlabel metal1 122 -817 231 -813 5 vdd
rlabel metal1 122 -907 231 -903 1 gnd
rlabel metal1 29 -840 29 -840 1 a3
rlabel metal1 27 -890 27 -890 1 b3
rlabel metal1 267 -866 267 -866 1 p3
rlabel metal1 173 -1128 173 -1128 1 gnd
rlabel metal1 185 -1052 185 -1052 5 vdd
rlabel metal1 118 -1093 118 -1093 1 a0
rlabel metal1 118 -1105 118 -1105 1 b0
rlabel metal1 174 -1215 174 -1215 1 gnd
rlabel metal1 186 -1139 186 -1139 5 vdd
rlabel metal1 119 -1180 119 -1180 1 a1
rlabel metal1 119 -1192 119 -1192 1 b1
rlabel metal1 176 -1303 176 -1303 1 gnd
rlabel metal1 188 -1227 188 -1227 5 vdd
rlabel metal1 121 -1268 121 -1268 1 a2
rlabel metal1 121 -1280 121 -1280 1 b2
rlabel metal1 176 -1389 176 -1389 1 gnd
rlabel metal1 188 -1313 188 -1313 5 vdd
rlabel metal1 121 -1354 121 -1354 1 a3
rlabel metal1 121 -1366 121 -1366 1 b3
rlabel metal1 635 -694 635 -694 1 gnd
rlabel metal1 647 -618 647 -618 5 vdd
rlabel metal1 580 -671 580 -671 1 c0
rlabel metal1 257 -1068 257 -1068 5 vdd!
rlabel metal1 263 -1113 263 -1113 1 gnd!
rlabel metal1 296 -1097 296 -1096 1 g0
rlabel metal1 257 -1155 257 -1155 5 vdd!
rlabel metal1 263 -1200 263 -1200 1 gnd!
rlabel metal1 260 -1243 260 -1243 5 vdd!
rlabel metal1 266 -1288 266 -1288 1 gnd!
rlabel metal1 261 -1329 261 -1329 5 vdd!
rlabel metal1 267 -1374 267 -1374 1 gnd!
rlabel metal1 299 -1272 299 -1272 1 g2
rlabel metal1 300 -1357 300 -1357 1 g3
rlabel metal1 723 -634 723 -634 5 vdd!
rlabel metal1 729 -679 729 -679 1 gnd!
rlabel metal1 796 -622 796 -622 5 vdd!
rlabel metal1 799 -687 799 -687 1 gnd!
rlabel metal1 833 -635 833 -635 5 vdd!
rlabel metal1 839 -680 839 -680 1 gnd!
rlabel metal1 887 -663 887 -663 1 c1
rlabel metal1 575 -782 575 -782 8 gnd
rlabel metal1 566 -705 566 -705 5 vdd
rlabel metal1 532 -752 533 -752 1 y
rlabel metal1 516 -703 517 -703 1 vdd
rlabel metal1 511 -793 512 -793 1 gnd
rlabel metal1 496 -885 496 -885 1 gnd
rlabel metal1 508 -809 508 -809 5 vdd
rlabel metal1 579 -825 579 -825 5 vdd!
rlabel metal1 585 -870 585 -870 1 gnd!
rlabel metal1 619 -742 619 -742 5 vdd!
rlabel metal1 622 -807 622 -807 1 gnd!
rlabel metal1 656 -755 656 -755 5 vdd!
rlabel metal1 662 -800 662 -800 1 gnd!
rlabel metal1 658 -850 658 -850 5 vdd!
rlabel metal1 661 -915 661 -915 1 gnd!
rlabel metal1 695 -863 695 -863 5 vdd!
rlabel metal1 701 -908 701 -908 1 gnd!
rlabel metal1 854 -1055 854 -1055 1 gnd
rlabel metal1 866 -979 866 -979 5 vdd
rlabel metal1 938 -995 938 -995 5 vdd!
rlabel metal1 944 -1040 944 -1040 1 gnd!
rlabel metal1 858 -1162 858 -1162 1 gnd
rlabel metal1 870 -1086 870 -1086 5 vdd
rlabel metal1 942 -1102 942 -1102 5 vdd!
rlabel metal1 948 -1147 948 -1147 1 gnd!
rlabel metal1 858 -1271 858 -1271 1 gnd
rlabel metal1 870 -1195 870 -1195 5 vdd
rlabel metal1 942 -1211 942 -1211 5 vdd!
rlabel metal1 948 -1256 948 -1256 1 gnd!
rlabel metal1 1018 -1045 1018 -1045 5 vdd!
rlabel metal1 1021 -1110 1021 -1110 1 gnd!
rlabel metal1 1055 -1058 1055 -1058 5 vdd!
rlabel metal1 1061 -1103 1061 -1103 1 gnd!
rlabel metal1 1018 -1214 1018 -1214 5 vdd!
rlabel metal1 1021 -1279 1021 -1279 1 gnd!
rlabel metal1 1055 -1227 1055 -1227 5 vdd!
rlabel metal1 1061 -1272 1061 -1272 1 gnd!
rlabel metal1 1106 -1124 1106 -1124 5 vdd!
rlabel metal1 1109 -1189 1109 -1189 1 gnd!
rlabel metal1 1143 -1137 1143 -1137 5 vdd!
rlabel metal1 1149 -1182 1149 -1182 1 gnd!
rlabel metal1 1186 -1166 1186 -1166 1 c3
rlabel metal1 1258 -1486 1258 -1486 1 gnd
rlabel metal1 1270 -1410 1270 -1410 5 vdd
rlabel metal1 1342 -1426 1342 -1426 5 vdd!
rlabel metal1 1348 -1471 1348 -1471 1 gnd!
rlabel metal1 1258 -1591 1258 -1591 1 gnd
rlabel metal1 1270 -1515 1270 -1515 5 vdd
rlabel metal1 1342 -1531 1342 -1531 5 vdd!
rlabel metal1 1348 -1576 1348 -1576 1 gnd!
rlabel metal1 1258 -1694 1258 -1694 1 gnd
rlabel metal1 1270 -1618 1270 -1618 5 vdd
rlabel metal1 1342 -1634 1342 -1634 5 vdd!
rlabel metal1 1348 -1679 1348 -1679 1 gnd!
rlabel metal1 1248 -1783 1248 -1783 1 gnd
rlabel metal1 1260 -1707 1260 -1707 5 vdd
rlabel metal1 1332 -1723 1332 -1723 5 vdd!
rlabel metal1 1338 -1768 1338 -1768 1 gnd!
rlabel metal1 1406 -1463 1406 -1463 5 vdd!
rlabel metal1 1409 -1528 1409 -1528 1 gnd!
rlabel metal1 1443 -1476 1443 -1476 5 vdd!
rlabel metal1 1449 -1521 1449 -1521 1 gnd!
rlabel metal1 1403 -1665 1403 -1665 5 vdd!
rlabel metal1 1406 -1730 1406 -1730 1 gnd!
rlabel metal1 1440 -1678 1440 -1678 5 vdd!
rlabel metal1 1446 -1723 1446 -1723 1 gnd!
rlabel metal1 1519 -1576 1519 -1576 5 vdd!
rlabel metal1 1522 -1641 1522 -1641 1 gnd!
rlabel metal1 1556 -1589 1556 -1589 5 vdd!
rlabel metal1 1562 -1634 1562 -1634 1 gnd!
rlabel metal1 1622 -1678 1622 -1678 5 vdd!
rlabel metal1 1625 -1743 1625 -1743 1 gnd!
rlabel metal1 1659 -1691 1659 -1691 5 vdd!
rlabel metal1 1665 -1736 1665 -1736 1 gnd!
rlabel metal1 1717 -1720 1717 -1720 1 c4
rlabel metal1 278 -1183 278 -1183 1 g1
rlabel metal1 225 -1357 225 -1357 1 test
rlabel metal1 711 -891 711 -891 1 c2
rlabel metal1 934 -525 1043 -521 5 vdd
rlabel metal1 934 -615 1043 -611 1 gnd
rlabel metal1 1103 -574 1103 -574 1 s0
rlabel metal1 944 -649 1053 -645 5 vdd
rlabel metal1 944 -739 1053 -735 1 gnd
rlabel metal1 1075 -697 1075 -697 1 s1
rlabel metal1 1292 -1089 1401 -1085 5 vdd
rlabel metal1 1292 -1179 1401 -1175 1 gnd
rlabel metal1 1434 -1138 1434 -1138 1 s3
rlabel metal1 848 -803 957 -799 5 vdd
rlabel metal1 848 -893 957 -889 1 gnd
rlabel metal1 980 -852 981 -851 1 s2
rlabel metal1 -344 -661 -344 -661 1 clk
rlabel metal1 -167 -482 -167 -482 5 vdd
rlabel metal1 -167 -647 -167 -647 1 gnd
rlabel metal1 -219 -482 -219 -482 5 vdd
rlabel metal1 -219 -647 -219 -647 1 gnd
rlabel metal1 -271 -647 -271 -647 1 gnd
rlabel metal1 -271 -482 -271 -482 5 vdd
rlabel metal1 -323 -647 -323 -647 1 gnd
rlabel metal1 -323 -482 -323 -482 5 vdd
rlabel metal1 -88 -630 -88 -630 1 gnd
rlabel metal1 -87 -528 -87 -528 5 vdd
rlabel metal1 -120 -630 -120 -630 1 gnd
rlabel metal1 -119 -528 -119 -528 5 vdd
rlabel metal1 -122 -757 -122 -757 5 vdd
rlabel metal1 -90 -757 -90 -757 5 vdd
rlabel metal1 -326 -711 -326 -711 5 vdd
rlabel metal1 -274 -711 -274 -711 5 vdd
rlabel metal1 -222 -711 -222 -711 5 vdd
rlabel metal1 -170 -711 -170 -711 5 vdd
rlabel metal1 -91 -859 -91 -859 1 gnd
rlabel metal1 -123 -859 -123 -859 1 gnd
rlabel metal1 -347 -890 -347 -890 1 clk
rlabel metal1 -170 -876 -170 -876 1 gnd
rlabel metal1 -222 -876 -222 -876 1 gnd
rlabel metal1 -274 -876 -274 -876 1 gnd
rlabel metal1 -326 -876 -326 -876 1 gnd
rlabel metal1 -347 -1106 -347 -1106 1 clk
rlabel metal1 -170 -927 -170 -927 5 vdd
rlabel metal1 -170 -1092 -170 -1092 1 gnd
rlabel metal1 -222 -927 -222 -927 5 vdd
rlabel metal1 -222 -1092 -222 -1092 1 gnd
rlabel metal1 -274 -1092 -274 -1092 1 gnd
rlabel metal1 -274 -927 -274 -927 5 vdd
rlabel metal1 -326 -1092 -326 -1092 1 gnd
rlabel metal1 -326 -927 -326 -927 5 vdd
rlabel metal1 -91 -1075 -91 -1075 1 gnd
rlabel metal1 -90 -973 -90 -973 5 vdd
rlabel metal1 -123 -1075 -123 -1075 1 gnd
rlabel metal1 -122 -973 -122 -973 5 vdd
rlabel metal1 -348 -1321 -348 -1321 1 clk
rlabel metal1 -171 -1142 -171 -1142 5 vdd
rlabel metal1 -171 -1307 -171 -1307 1 gnd
rlabel metal1 -223 -1142 -223 -1142 5 vdd
rlabel metal1 -223 -1307 -223 -1307 1 gnd
rlabel metal1 -275 -1307 -275 -1307 1 gnd
rlabel metal1 -275 -1142 -275 -1142 5 vdd
rlabel metal1 -327 -1307 -327 -1307 1 gnd
rlabel metal1 -327 -1142 -327 -1142 5 vdd
rlabel metal1 -92 -1290 -92 -1290 1 gnd
rlabel metal1 -91 -1188 -91 -1188 5 vdd
rlabel metal1 -124 -1290 -124 -1290 1 gnd
rlabel metal1 -123 -1188 -123 -1188 5 vdd
rlabel metal1 -356 -1551 -356 -1551 1 clk
rlabel metal1 -179 -1372 -179 -1372 5 vdd
rlabel metal1 -179 -1537 -179 -1537 1 gnd
rlabel metal1 -231 -1372 -231 -1372 5 vdd
rlabel metal1 -231 -1537 -231 -1537 1 gnd
rlabel metal1 -283 -1537 -283 -1537 1 gnd
rlabel metal1 -283 -1372 -283 -1372 5 vdd
rlabel metal1 -335 -1537 -335 -1537 1 gnd
rlabel metal1 -335 -1372 -335 -1372 5 vdd
rlabel metal1 -100 -1520 -100 -1520 1 gnd
rlabel metal1 -99 -1418 -99 -1418 5 vdd
rlabel metal1 -132 -1520 -132 -1520 1 gnd
rlabel metal1 -131 -1418 -131 -1418 5 vdd
rlabel metal1 -354 -1777 -354 -1777 1 clk
rlabel metal1 -177 -1598 -177 -1598 5 vdd
rlabel metal1 -177 -1763 -177 -1763 1 gnd
rlabel metal1 -229 -1598 -229 -1598 5 vdd
rlabel metal1 -229 -1763 -229 -1763 1 gnd
rlabel metal1 -281 -1763 -281 -1763 1 gnd
rlabel metal1 -281 -1598 -281 -1598 5 vdd
rlabel metal1 -333 -1763 -333 -1763 1 gnd
rlabel metal1 -333 -1598 -333 -1598 5 vdd
rlabel metal1 -98 -1746 -98 -1746 1 gnd
rlabel metal1 -97 -1644 -97 -1644 5 vdd
rlabel metal1 -130 -1746 -130 -1746 1 gnd
rlabel metal1 -129 -1644 -129 -1644 5 vdd
rlabel metal1 -354 -2000 -354 -2000 1 clk
rlabel metal1 -177 -1821 -177 -1821 5 vdd
rlabel metal1 -177 -1986 -177 -1986 1 gnd
rlabel metal1 -229 -1821 -229 -1821 5 vdd
rlabel metal1 -229 -1986 -229 -1986 1 gnd
rlabel metal1 -281 -1986 -281 -1986 1 gnd
rlabel metal1 -281 -1821 -281 -1821 5 vdd
rlabel metal1 -333 -1986 -333 -1986 1 gnd
rlabel metal1 -333 -1821 -333 -1821 5 vdd
rlabel metal1 -98 -1969 -98 -1969 1 gnd
rlabel metal1 -97 -1867 -97 -1867 5 vdd
rlabel metal1 -130 -1969 -130 -1969 1 gnd
rlabel metal1 -129 -1867 -129 -1867 5 vdd
rlabel metal1 -341 -434 -341 -434 1 clk
rlabel metal1 -164 -255 -164 -255 5 vdd
rlabel metal1 -164 -420 -164 -420 1 gnd
rlabel metal1 -216 -255 -216 -255 5 vdd
rlabel metal1 -216 -420 -216 -420 1 gnd
rlabel metal1 -268 -420 -268 -420 1 gnd
rlabel metal1 -268 -255 -268 -255 5 vdd
rlabel metal1 -320 -420 -320 -420 1 gnd
rlabel metal1 -320 -255 -320 -255 5 vdd
rlabel metal1 -85 -403 -85 -403 1 gnd
rlabel metal1 -84 -301 -84 -301 5 vdd
rlabel metal1 -117 -403 -117 -403 1 gnd
rlabel metal1 -116 -301 -116 -301 5 vdd
rlabel metal1 -358 -347 -358 -347 1 a00
rlabel metal1 -55 -366 -55 -366 1 a0
rlabel metal1 -363 -573 -363 -573 1 a11
rlabel metal1 -59 -594 -59 -594 1 a1
rlabel metal1 -364 -803 -364 -803 1 a22
rlabel metal1 -63 -822 -63 -822 1 a2
rlabel metal1 -364 -1018 -364 -1018 1 a33
rlabel metal1 -61 -1038 -61 -1038 1 a3
rlabel metal1 -366 -1233 -366 -1233 1 b00
rlabel metal1 -63 -1254 -63 -1254 1 b0
rlabel metal1 -373 -1463 -373 -1463 3 b11
rlabel metal1 -70 -1484 -70 -1484 1 b1
rlabel metal1 -370 -1688 -370 -1688 1 b22
rlabel metal1 -69 -1710 -69 -1710 1 b2
rlabel metal1 -371 -1912 -371 -1912 1 b33
rlabel metal1 -69 -1933 -69 -1933 1 b3
rlabel metal1 1559 -926 1559 -926 1 clk
rlabel metal1 1736 -747 1736 -747 5 vdd
rlabel metal1 1736 -912 1736 -912 1 gnd
rlabel metal1 1684 -747 1684 -747 5 vdd
rlabel metal1 1684 -912 1684 -912 1 gnd
rlabel metal1 1632 -912 1632 -912 1 gnd
rlabel metal1 1632 -747 1632 -747 5 vdd
rlabel metal1 1580 -912 1580 -912 1 gnd
rlabel metal1 1580 -747 1580 -747 5 vdd
rlabel metal1 1815 -895 1815 -895 1 gnd
rlabel metal1 1816 -793 1816 -793 5 vdd
rlabel metal1 1783 -895 1783 -895 1 gnd
rlabel metal1 1784 -793 1784 -793 5 vdd
rlabel metal1 1559 -1159 1559 -1159 1 clk
rlabel metal1 1736 -980 1736 -980 5 vdd
rlabel metal1 1736 -1145 1736 -1145 1 gnd
rlabel metal1 1684 -980 1684 -980 5 vdd
rlabel metal1 1684 -1145 1684 -1145 1 gnd
rlabel metal1 1632 -1145 1632 -1145 1 gnd
rlabel metal1 1632 -980 1632 -980 5 vdd
rlabel metal1 1580 -1145 1580 -1145 1 gnd
rlabel metal1 1580 -980 1580 -980 5 vdd
rlabel metal1 1815 -1128 1815 -1128 1 gnd
rlabel metal1 1816 -1026 1816 -1026 5 vdd
rlabel metal1 1783 -1128 1783 -1128 1 gnd
rlabel metal1 1784 -1026 1784 -1026 5 vdd
rlabel metal1 1554 -1385 1554 -1385 1 clk
rlabel metal1 1731 -1206 1731 -1206 5 vdd
rlabel metal1 1731 -1371 1731 -1371 1 gnd
rlabel metal1 1679 -1206 1679 -1206 5 vdd
rlabel metal1 1679 -1371 1679 -1371 1 gnd
rlabel metal1 1627 -1371 1627 -1371 1 gnd
rlabel metal1 1627 -1206 1627 -1206 5 vdd
rlabel metal1 1575 -1371 1575 -1371 1 gnd
rlabel metal1 1575 -1206 1575 -1206 5 vdd
rlabel metal1 1810 -1354 1810 -1354 1 gnd
rlabel metal1 1811 -1252 1811 -1252 5 vdd
rlabel metal1 1778 -1354 1778 -1354 1 gnd
rlabel metal1 1779 -1252 1779 -1252 5 vdd
rlabel metal1 1566 -448 1566 -448 1 clk
rlabel metal1 1743 -269 1743 -269 5 vdd
rlabel metal1 1743 -434 1743 -434 1 gnd
rlabel metal1 1691 -269 1691 -269 5 vdd
rlabel metal1 1691 -434 1691 -434 1 gnd
rlabel metal1 1639 -434 1639 -434 1 gnd
rlabel metal1 1639 -269 1639 -269 5 vdd
rlabel metal1 1587 -434 1587 -434 1 gnd
rlabel metal1 1587 -269 1587 -269 5 vdd
rlabel metal1 1822 -417 1822 -417 1 gnd
rlabel metal1 1823 -315 1823 -315 5 vdd
rlabel metal1 1790 -417 1790 -417 1 gnd
rlabel metal1 1791 -315 1791 -315 5 vdd
rlabel metal1 1558 -690 1558 -690 1 clk
rlabel metal1 1735 -511 1735 -511 5 vdd
rlabel metal1 1735 -676 1735 -676 1 gnd
rlabel metal1 1683 -511 1683 -511 5 vdd
rlabel metal1 1683 -676 1683 -676 1 gnd
rlabel metal1 1631 -676 1631 -676 1 gnd
rlabel metal1 1631 -511 1631 -511 5 vdd
rlabel metal1 1579 -676 1579 -676 1 gnd
rlabel metal1 1579 -511 1579 -511 5 vdd
rlabel metal1 1814 -659 1814 -659 1 gnd
rlabel metal1 1815 -557 1815 -557 5 vdd
rlabel metal1 1782 -659 1782 -659 1 gnd
rlabel metal1 1783 -557 1783 -557 5 vdd
rlabel metal1 1852 -380 1852 -380 1 s00
rlabel metal1 1550 -361 1550 -361 1 s0
rlabel metal1 1844 -622 1844 -622 1 s11
rlabel metal1 1544 -603 1544 -603 1 s1
rlabel metal1 1844 -858 1844 -858 1 s22
rlabel metal1 1543 -838 1543 -838 1 s2
rlabel metal1 1843 -1092 1843 -1092 1 s33
rlabel metal1 1542 -1071 1542 -1071 1 s3
rlabel metal1 1839 -1317 1839 -1317 1 c44
rlabel metal1 1539 -1297 1539 -1297 1 c4
<< end >>
