magic
tech scmos
timestamp 1731850112
<< nwell >>
rect 0 0 40 34
<< ntransistor >>
rect 12 -38 15 -22
rect 25 -38 28 -22
<< ptransistor >>
rect 12 6 15 26
rect 25 6 28 26
<< ndiffusion >>
rect 10 -27 12 -22
rect 6 -38 12 -27
rect 15 -38 25 -22
rect 28 -27 30 -22
rect 28 -38 34 -27
<< pdiffusion >>
rect 10 21 12 26
rect 6 6 12 21
rect 15 21 18 26
rect 22 21 25 26
rect 15 6 25 21
rect 28 21 30 26
rect 28 6 34 21
<< ndcontact >>
rect 6 -27 10 -22
rect 30 -27 34 -22
<< pdcontact >>
rect 6 21 10 26
rect 18 21 22 26
rect 30 21 34 26
<< polysilicon >>
rect 12 26 15 30
rect 25 26 28 30
rect 12 -3 15 6
rect 14 -7 15 -3
rect 12 -22 15 -7
rect 25 -14 28 6
rect 27 -18 28 -14
rect 25 -22 28 -18
rect 12 -43 15 -38
rect 25 -43 28 -38
<< polycontact >>
rect 10 -7 14 -3
rect 22 -18 27 -14
<< metal1 >>
rect 6 34 34 38
rect 6 26 10 34
rect 30 26 34 34
rect 6 -7 10 -3
rect 18 -7 22 21
rect 18 -11 34 -7
rect 6 -18 22 -14
rect 27 -18 28 -14
rect 6 -19 28 -18
rect 31 -22 34 -11
rect 6 -42 10 -27
<< labels >>
rlabel metal1 7 -5 7 -5 1 a
rlabel metal1 8 -16 8 -16 1 b
rlabel metal1 33 -9 33 -9 1 out
rlabel metal1 8 -40 8 -40 1 gnd
rlabel metal1 20 36 20 36 5 vdd
<< end >>
