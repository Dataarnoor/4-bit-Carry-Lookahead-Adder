magic
tech scmos
timestamp 1732046546
<< nwell >>
rect 439 69 471 195
rect 491 69 523 195
rect 543 131 575 195
rect 595 131 627 195
rect 648 86 712 150
<< ntransistor >>
rect 558 84 560 104
rect 610 84 612 104
rect 454 37 456 57
rect 506 37 508 57
rect 558 37 560 57
rect 610 37 612 57
rect 663 55 665 75
rect 695 55 697 75
<< ptransistor >>
rect 454 140 456 180
rect 506 140 508 180
rect 558 140 560 180
rect 610 140 612 180
rect 454 78 456 118
rect 506 78 508 118
rect 663 95 665 135
rect 695 95 697 135
<< ndiffusion >>
rect 557 84 558 104
rect 560 84 561 104
rect 609 84 610 104
rect 612 84 613 104
rect 453 37 454 57
rect 456 37 457 57
rect 505 37 506 57
rect 508 37 509 57
rect 557 37 558 57
rect 560 37 561 57
rect 609 37 610 57
rect 612 37 613 57
rect 662 55 663 75
rect 665 55 666 75
rect 694 55 695 75
rect 697 55 698 75
<< pdiffusion >>
rect 453 140 454 180
rect 456 140 457 180
rect 505 140 506 180
rect 508 140 509 180
rect 557 140 558 180
rect 560 140 561 180
rect 609 140 610 180
rect 612 140 613 180
rect 453 78 454 118
rect 456 78 457 118
rect 505 78 506 118
rect 508 78 509 118
rect 662 95 663 135
rect 665 95 666 135
rect 694 95 695 135
rect 697 95 698 135
<< ndcontact >>
rect 553 84 557 104
rect 561 84 565 104
rect 605 84 609 104
rect 613 84 617 104
rect 449 37 453 57
rect 457 37 461 57
rect 501 37 505 57
rect 509 37 513 57
rect 553 37 557 57
rect 561 37 565 57
rect 605 37 609 57
rect 613 37 617 57
rect 658 55 662 75
rect 666 55 670 75
rect 690 55 694 75
rect 698 55 702 75
<< pdcontact >>
rect 449 140 453 180
rect 457 140 461 180
rect 501 140 505 180
rect 509 140 513 180
rect 553 140 557 180
rect 561 140 565 180
rect 605 140 609 180
rect 613 140 617 180
rect 449 78 453 118
rect 457 78 461 118
rect 501 78 505 118
rect 509 78 513 118
rect 658 95 662 135
rect 666 95 670 135
rect 690 95 694 135
rect 698 95 702 135
<< psubstratepcontact >>
rect 650 42 654 46
rect 674 42 678 46
rect 682 42 686 46
rect 706 42 710 46
rect 466 24 470 28
rect 518 24 522 28
rect 570 24 574 28
rect 622 24 626 28
<< nsubstratencontact >>
rect 442 188 446 192
rect 464 188 468 192
rect 494 188 498 192
rect 516 188 520 192
rect 546 188 550 192
rect 568 188 572 192
rect 598 188 602 192
rect 620 188 624 192
rect 651 143 655 147
rect 673 143 677 147
rect 683 143 687 147
rect 705 143 709 147
<< polysilicon >>
rect 454 180 456 184
rect 506 180 508 184
rect 558 180 560 184
rect 610 180 612 184
rect 454 131 456 140
rect 506 131 508 140
rect 558 131 560 140
rect 610 131 612 140
rect 663 135 665 139
rect 695 135 697 139
rect 454 118 456 122
rect 506 118 508 122
rect 558 104 560 113
rect 610 104 612 113
rect 558 81 560 84
rect 610 81 612 84
rect 454 69 456 78
rect 506 69 508 78
rect 663 75 665 95
rect 695 75 697 95
rect 454 57 456 65
rect 506 57 508 65
rect 558 57 560 65
rect 610 57 612 65
rect 663 51 665 55
rect 695 51 697 55
rect 454 33 456 37
rect 506 33 508 37
rect 558 33 560 37
rect 610 33 612 37
<< polycontact >>
rect 449 131 454 136
rect 501 131 506 136
rect 553 131 558 136
rect 605 131 610 136
rect 553 108 558 113
rect 605 108 610 113
rect 658 78 663 83
rect 449 69 454 74
rect 501 69 506 74
rect 690 78 695 83
rect 449 60 454 65
rect 501 60 506 65
rect 553 60 558 65
rect 605 60 610 65
<< metal1 >>
rect 439 192 627 195
rect 439 188 442 192
rect 446 188 464 192
rect 468 188 494 192
rect 498 188 516 192
rect 520 188 546 192
rect 550 188 568 192
rect 572 188 598 192
rect 602 188 620 192
rect 624 188 627 192
rect 439 186 627 188
rect 449 180 453 186
rect 501 180 505 186
rect 553 180 557 186
rect 605 180 609 186
rect 648 147 712 150
rect 648 143 651 147
rect 655 143 673 147
rect 677 143 683 147
rect 687 143 705 147
rect 709 143 712 147
rect 648 141 712 143
rect 426 131 449 136
rect 426 65 431 131
rect 457 127 461 140
rect 449 123 461 127
rect 479 131 501 136
rect 449 118 453 123
rect 444 69 449 74
rect 457 65 461 78
rect 479 65 484 131
rect 509 127 513 140
rect 561 136 565 140
rect 613 136 617 140
rect 501 123 513 127
rect 531 131 553 136
rect 561 131 605 136
rect 613 131 637 136
rect 501 118 505 123
rect 496 69 501 74
rect 509 65 513 78
rect 531 65 536 131
rect 550 108 553 113
rect 561 104 565 131
rect 553 73 557 84
rect 553 69 565 73
rect 426 60 449 65
rect 457 60 501 65
rect 509 60 553 65
rect 457 57 461 60
rect 509 57 513 60
rect 561 57 565 69
rect 583 65 588 131
rect 602 108 605 113
rect 613 104 617 131
rect 605 73 609 84
rect 632 83 637 131
rect 658 135 662 141
rect 690 135 694 141
rect 666 83 670 95
rect 698 83 702 95
rect 632 78 658 83
rect 666 78 690 83
rect 698 78 712 83
rect 666 75 670 78
rect 698 75 702 78
rect 605 69 617 73
rect 583 60 605 65
rect 613 57 617 69
rect 658 48 662 55
rect 690 48 694 55
rect 648 46 712 48
rect 648 42 650 46
rect 654 42 674 46
rect 678 42 682 46
rect 686 42 706 46
rect 710 42 712 46
rect 648 40 712 42
rect 449 29 453 37
rect 501 29 505 37
rect 553 29 557 37
rect 605 29 609 37
rect 439 28 627 29
rect 439 24 466 28
rect 470 24 518 28
rect 522 24 570 28
rect 574 24 622 28
rect 626 24 627 28
rect 439 23 627 24
rect 432 10 439 15
rect 444 10 491 15
rect 496 10 545 15
rect 550 10 597 15
<< m2contact >>
rect 439 69 444 74
rect 491 69 496 74
rect 545 108 550 113
rect 597 108 602 113
rect 439 10 444 15
rect 491 10 496 15
rect 545 10 550 15
rect 597 10 602 15
<< metal2 >>
rect 439 15 444 69
rect 491 15 496 69
rect 545 15 550 108
rect 597 15 602 108
<< labels >>
rlabel metal1 455 191 455 191 5 vdd
rlabel metal1 455 26 455 26 1 gnd
rlabel metal1 507 191 507 191 5 vdd
rlabel metal1 507 26 507 26 1 gnd
rlabel metal1 559 26 559 26 1 gnd
rlabel metal1 559 191 559 191 5 vdd
rlabel metal1 611 26 611 26 1 gnd
rlabel metal1 611 191 611 191 5 vdd
rlabel metal1 428 101 428 101 1 d
rlabel metal1 434 12 434 12 1 clk
rlabel metal1 695 44 695 44 1 gnd
rlabel metal1 696 146 696 146 5 vdd
rlabel metal1 663 44 663 44 1 gnd
rlabel metal1 664 146 664 146 5 vdd
rlabel metal1 708 81 708 81 7 q
<< end >>
